* SPICE3 file created from XNOR.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'




.option scale=1u

M1000 a_n100_18# Vb Vdd w_n115_16# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1001 Vdd a_n100_18# a_n33_n26# w_n48_n28# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1002 a_35_22# a_n33_n26# Vdd w_20_20# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1003 Vdd a_n33_57# a_35_22# w_20_20# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1004 a_35_22# a_n33_57# a_35_n18# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1005 a_n33_57# a_n100_18# Vdd w_n48_55# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1006 Vdd Va a_n33_57# w_n48_55# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1007 a_n100_18# Va a_n100_n22# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1008 a_n100_n22# Vb gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1009 a_n33_n66# Vb gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1010 a_n33_17# a_n100_18# gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1011 a_n33_57# Va a_n33_17# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1012 Vout a_35_22# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1013 a_35_n18# a_n33_n26# gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1014 Vout a_35_22# Vdd w_93_11# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1015 a_n33_n26# Vb Vdd w_n48_n28# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1016 Vdd Va a_n100_18# w_n115_16# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1017 a_n33_n26# a_n100_18# a_n33_n66# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
C0 Vout 0 3.76f 
C1 a_35_22# 0 22.652f 
C2 gnd 0 70.304f 
C3 a_n33_n26# 0 35.45f 
C4 Vb 0 55.483997f 
C5 a_n33_57# 0 36.766f 
C6 Va 0 60.888996f 
C7 a_n100_18# 0 60.184002f 
C8 Vdd 0 61.128002f 

Va Va gnd 1
Vb Vb gnd 0


.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(Va) v(Vb)+2 v(Vout)+4 
.end
.endc