Decoder Implementation

.include TSMC_180nm.txt
.include NAND.sub
.include NOT.sub
.include AND.sub
.include 3AND.sub
.include 4AND.sub
.include 5AND.sub
.include OR.sub
.include 3OR.sub
.include 4OR.sub
.include XOR.sub
.include XNOR.sub
.include FullAdder.sub
.include Adder.sub
.include Sub.sub
.include Comparator.sub
.include ENABLE.sub
.include ANDING.sub
.include DECODER.sub


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_c c gnd dc 0
V_in_cin1 cin1 gnd dc 0
V_in_cin0 cin0 gnd dc 1.8
V_in_s0 s0 gnd dc 1.8
V_in_s1 s1 gnd dc 0

V_in_a3 a3 gnd dc 1.8
V_in_a2 a2 gnd dc 1.8
V_in_a1 a1 gnd dc 1.8
V_in_a0 a0 gnd dc 0


V_in_b3 b3 gnd dc 0
V_in_b2 b2 gnd dc 1.8
V_in_b1 b1 gnd dc 1.8
V_in_b0 b0 gnd dc 1.8



X1 a3 a2 a1 a0 b3 b2 b1 b0 s1 s0 c y03 y02 y01 y00 cout cin0 cin1 y13 y12 y11 y10 si ga gb e y33 y32 y31 y30 node_x gnd DECODER

.tran 1n 800n

.control
run


* plot v(cout)+2 v(si)+4
* plot v(a3) v(b3)+2 v(y03)+4 v(y13)+6 v(y33)+8
* plot v(a2) v(b2)+2 v(y02)+4 v(y12)+6 v(y32)+8
* plot v(a1) v(b1)+2 v(y01)+4 v(y11)+6 v(y31)+8
* plot v(a0) v(b0)+2 v(y00)+4 v(y10)+6 v(y30)+8
* plot v(ga) v(gb)+2 v(e)+4

plot v(y10) v(y11)+2 v(y12)+4 v(y13)+6 v(si)+8

.end
.endc
