* SPICE3 file created from NOTANDGATE.ext - technology: scmos


.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'


.option scale=1u

M1000 Vout a_15_50# Vdd w_n26_48# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1001 a_n12_10# Vb gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1002 Vout a_15_50# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1003 a_15_50# a_n12_10# Vdd w_n26_48# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1004 Vdd Va a_15_50# w_n26_48# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1005 a_15_10# a_n12_10# gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1006 a_15_50# Va a_15_10# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1007 a_n12_10# Vb Vdd w_n26_48# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
C0 gnd 0 16.168001f 
C1 Vout 0 6.392f 
C2 a_15_50# 0 21.108f 
C3 Va 0 20.682f 
C4 a_n12_10# 0 20.786001f 
C5 Vb 0 12.46f 
C6 Vdd 0 17.672f 



Va Va gnd 1
Vb Vb gnd 0


.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(Va) v(Vb)+2 v(Vout)+4 
.end
.endc