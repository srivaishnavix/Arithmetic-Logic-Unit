magic
tech scmos
timestamp 1701017107
<< nwell >>
rect -476 132 -434 144
rect -241 132 -199 144
rect 47 132 89 144
rect 282 132 324 144
rect 570 132 612 144
rect 805 132 847 144
rect 1093 132 1135 144
rect 1328 132 1370 144
rect -543 93 -501 105
rect -408 97 -366 109
rect -308 93 -266 105
rect -173 97 -131 109
rect -20 93 22 105
rect 115 97 157 109
rect 215 93 257 105
rect 350 97 392 109
rect 503 93 545 105
rect 638 97 680 109
rect 738 93 780 105
rect 873 97 915 109
rect 1026 93 1068 105
rect 1161 97 1203 109
rect 1261 93 1303 105
rect 1396 97 1438 109
rect -476 49 -434 61
rect -241 49 -199 61
rect 47 49 89 61
rect 282 49 324 61
rect 570 49 612 61
rect 805 49 847 61
rect 1093 49 1135 61
rect 1328 49 1370 61
rect -562 -41 -494 -29
rect -310 -41 -242 -29
rect -193 -41 -125 -29
rect -39 -41 29 -29
rect 213 -41 281 -29
rect 330 -41 398 -29
rect 484 -41 552 -29
rect 736 -41 804 -29
rect 853 -41 921 -29
rect 1007 -41 1075 -29
rect 1259 -41 1327 -29
rect 1376 -41 1444 -29
<< polysilicon >>
rect -598 74 -594 165
rect -590 82 -586 165
rect -464 142 -461 146
rect -449 142 -446 146
rect -229 142 -226 146
rect -214 142 -211 146
rect -464 111 -461 134
rect -449 119 -446 134
rect -450 115 -446 119
rect -465 107 -461 111
rect -531 103 -528 107
rect -516 103 -513 107
rect -464 102 -461 107
rect -449 102 -446 115
rect -229 111 -226 134
rect -214 119 -211 134
rect -215 115 -211 119
rect -396 107 -393 111
rect -381 107 -378 111
rect -230 107 -226 111
rect -572 86 -561 89
rect -572 -25 -569 86
rect -564 83 -561 86
rect -564 82 -560 83
rect -531 72 -528 95
rect -516 80 -513 95
rect -296 103 -293 107
rect -281 103 -278 107
rect -464 92 -461 94
rect -449 92 -446 94
rect -517 76 -513 80
rect -396 76 -393 99
rect -381 84 -378 99
rect -229 102 -226 107
rect -214 102 -211 115
rect -161 107 -158 111
rect -146 107 -143 111
rect -382 80 -378 84
rect -532 68 -528 72
rect -564 65 -560 66
rect -564 23 -561 65
rect -531 63 -528 68
rect -516 63 -513 76
rect -397 72 -393 76
rect -396 67 -393 72
rect -381 67 -378 80
rect -464 59 -461 63
rect -449 59 -446 63
rect -531 53 -528 55
rect -516 53 -513 55
rect -396 57 -393 59
rect -381 57 -378 59
rect -464 28 -461 51
rect -449 36 -446 51
rect -450 32 -446 36
rect -465 24 -461 28
rect -564 20 -539 23
rect -542 -25 -539 20
rect -464 19 -461 24
rect -449 19 -446 32
rect -464 9 -461 11
rect -449 9 -446 11
rect -572 -28 -547 -25
rect -542 -28 -532 -25
rect -550 -31 -547 -28
rect -535 -31 -532 -28
rect -508 -31 -506 -27
rect -550 -71 -547 -39
rect -535 -71 -532 -39
rect -508 -71 -506 -39
rect -550 -81 -547 -79
rect -535 -81 -532 -79
rect -508 -81 -506 -79
rect -492 -93 -488 -52
rect -357 -62 -353 -13
rect -345 -46 -341 78
rect -296 72 -293 95
rect -281 80 -278 95
rect -229 92 -226 94
rect -214 92 -211 94
rect -282 76 -278 80
rect -161 76 -158 99
rect -146 84 -143 99
rect -147 80 -143 84
rect -297 68 -293 72
rect -331 -5 -327 66
rect -296 63 -293 68
rect -281 63 -278 76
rect -162 72 -158 76
rect -161 67 -158 72
rect -146 67 -143 80
rect -229 59 -226 63
rect -214 59 -211 63
rect -296 53 -293 55
rect -281 53 -278 55
rect -161 57 -158 59
rect -146 57 -143 59
rect -229 28 -226 51
rect -214 36 -211 51
rect -215 32 -211 36
rect -230 24 -226 28
rect -229 19 -226 24
rect -214 19 -211 32
rect -229 9 -226 11
rect -214 9 -211 11
rect -298 -31 -295 -27
rect -283 -31 -280 -27
rect -256 -31 -254 -27
rect -181 -31 -178 -27
rect -166 -31 -163 -27
rect -139 -31 -137 -27
rect -345 -50 -343 -46
rect -298 -62 -295 -39
rect -283 -54 -280 -39
rect -284 -58 -280 -54
rect -357 -66 -355 -62
rect -299 -66 -295 -62
rect -298 -71 -295 -66
rect -283 -71 -280 -58
rect -256 -71 -254 -39
rect -181 -62 -178 -39
rect -182 -66 -178 -62
rect -181 -71 -178 -66
rect -166 -71 -163 -39
rect -139 -71 -137 -39
rect -298 -81 -295 -79
rect -283 -81 -280 -79
rect -256 -81 -254 -79
rect -181 -81 -178 -79
rect -166 -81 -163 -79
rect -139 -81 -137 -79
rect -181 -83 -174 -81
rect -177 -93 -174 -83
rect -492 -97 -174 -93
rect -104 -104 -100 78
rect -75 74 -71 165
rect -67 82 -63 165
rect 59 142 62 146
rect 74 142 77 146
rect 294 142 297 146
rect 309 142 312 146
rect 59 111 62 134
rect 74 119 77 134
rect 73 115 77 119
rect 58 107 62 111
rect -8 103 -5 107
rect 7 103 10 107
rect 59 102 62 107
rect 74 102 77 115
rect 294 111 297 134
rect 309 119 312 134
rect 308 115 312 119
rect 127 107 130 111
rect 142 107 145 111
rect 293 107 297 111
rect -49 86 -38 89
rect -49 -25 -46 86
rect -41 83 -38 86
rect -41 82 -37 83
rect -8 72 -5 95
rect 7 80 10 95
rect 227 103 230 107
rect 242 103 245 107
rect 59 92 62 94
rect 74 92 77 94
rect 6 76 10 80
rect 127 76 130 99
rect 142 84 145 99
rect 294 102 297 107
rect 309 102 312 115
rect 362 107 365 111
rect 377 107 380 111
rect 141 80 145 84
rect -9 68 -5 72
rect -41 65 -37 66
rect -41 23 -38 65
rect -8 63 -5 68
rect 7 63 10 76
rect 126 72 130 76
rect 127 67 130 72
rect 142 67 145 80
rect 59 59 62 63
rect 74 59 77 63
rect -8 53 -5 55
rect 7 53 10 55
rect 127 57 130 59
rect 142 57 145 59
rect 59 28 62 51
rect 74 36 77 51
rect 73 32 77 36
rect 58 24 62 28
rect -41 20 -16 23
rect -19 -25 -16 20
rect 59 19 62 24
rect 74 19 77 32
rect 59 9 62 11
rect 74 9 77 11
rect -49 -28 -24 -25
rect -19 -28 -9 -25
rect -27 -31 -24 -28
rect -12 -31 -9 -28
rect 15 -31 17 -27
rect -27 -71 -24 -39
rect -12 -71 -9 -39
rect 15 -71 17 -39
rect -27 -81 -24 -79
rect -12 -81 -9 -79
rect 15 -81 17 -79
rect 31 -93 35 -52
rect 166 -62 170 -13
rect 178 -46 182 78
rect 227 72 230 95
rect 242 80 245 95
rect 294 92 297 94
rect 309 92 312 94
rect 241 76 245 80
rect 362 76 365 99
rect 377 84 380 99
rect 376 80 380 84
rect 226 68 230 72
rect 192 -5 196 66
rect 227 63 230 68
rect 242 63 245 76
rect 361 72 365 76
rect 362 67 365 72
rect 377 67 380 80
rect 294 59 297 63
rect 309 59 312 63
rect 227 53 230 55
rect 242 53 245 55
rect 362 57 365 59
rect 377 57 380 59
rect 294 28 297 51
rect 309 36 312 51
rect 308 32 312 36
rect 293 24 297 28
rect 294 19 297 24
rect 309 19 312 32
rect 294 9 297 11
rect 309 9 312 11
rect 225 -31 228 -27
rect 240 -31 243 -27
rect 267 -31 269 -27
rect 342 -31 345 -27
rect 357 -31 360 -27
rect 384 -31 386 -27
rect 178 -50 180 -46
rect 225 -62 228 -39
rect 240 -54 243 -39
rect 239 -58 243 -54
rect 166 -66 168 -62
rect 224 -66 228 -62
rect 225 -71 228 -66
rect 240 -71 243 -58
rect 267 -71 269 -39
rect 342 -62 345 -39
rect 341 -66 345 -62
rect 342 -71 345 -66
rect 357 -71 360 -39
rect 384 -71 386 -39
rect 225 -81 228 -79
rect 240 -81 243 -79
rect 267 -81 269 -79
rect 342 -81 345 -79
rect 357 -81 360 -79
rect 384 -81 386 -79
rect 342 -83 349 -81
rect 346 -93 349 -83
rect 31 -97 349 -93
rect 419 -104 423 78
rect 448 74 452 165
rect 456 82 460 165
rect 582 142 585 146
rect 597 142 600 146
rect 817 142 820 146
rect 832 142 835 146
rect 582 111 585 134
rect 597 119 600 134
rect 596 115 600 119
rect 581 107 585 111
rect 515 103 518 107
rect 530 103 533 107
rect 582 102 585 107
rect 597 102 600 115
rect 817 111 820 134
rect 832 119 835 134
rect 831 115 835 119
rect 650 107 653 111
rect 665 107 668 111
rect 816 107 820 111
rect 474 86 485 89
rect 474 -25 477 86
rect 482 83 485 86
rect 482 82 486 83
rect 515 72 518 95
rect 530 80 533 95
rect 750 103 753 107
rect 765 103 768 107
rect 582 92 585 94
rect 597 92 600 94
rect 529 76 533 80
rect 650 76 653 99
rect 665 84 668 99
rect 817 102 820 107
rect 832 102 835 115
rect 885 107 888 111
rect 900 107 903 111
rect 664 80 668 84
rect 514 68 518 72
rect 482 65 486 66
rect 482 23 485 65
rect 515 63 518 68
rect 530 63 533 76
rect 649 72 653 76
rect 650 67 653 72
rect 665 67 668 80
rect 582 59 585 63
rect 597 59 600 63
rect 515 53 518 55
rect 530 53 533 55
rect 650 57 653 59
rect 665 57 668 59
rect 582 28 585 51
rect 597 36 600 51
rect 596 32 600 36
rect 581 24 585 28
rect 482 20 507 23
rect 504 -25 507 20
rect 582 19 585 24
rect 597 19 600 32
rect 582 9 585 11
rect 597 9 600 11
rect 474 -28 499 -25
rect 504 -28 514 -25
rect 496 -31 499 -28
rect 511 -31 514 -28
rect 538 -31 540 -27
rect 496 -71 499 -39
rect 511 -71 514 -39
rect 538 -71 540 -39
rect 496 -81 499 -79
rect 511 -81 514 -79
rect 538 -81 540 -79
rect 554 -93 558 -52
rect 689 -62 693 -13
rect 701 -46 705 78
rect 750 72 753 95
rect 765 80 768 95
rect 817 92 820 94
rect 832 92 835 94
rect 764 76 768 80
rect 885 76 888 99
rect 900 84 903 99
rect 899 80 903 84
rect 749 68 753 72
rect 715 -5 719 66
rect 750 63 753 68
rect 765 63 768 76
rect 884 72 888 76
rect 885 67 888 72
rect 900 67 903 80
rect 817 59 820 63
rect 832 59 835 63
rect 750 53 753 55
rect 765 53 768 55
rect 885 57 888 59
rect 900 57 903 59
rect 817 28 820 51
rect 832 36 835 51
rect 831 32 835 36
rect 816 24 820 28
rect 817 19 820 24
rect 832 19 835 32
rect 817 9 820 11
rect 832 9 835 11
rect 748 -31 751 -27
rect 763 -31 766 -27
rect 790 -31 792 -27
rect 865 -31 868 -27
rect 880 -31 883 -27
rect 907 -31 909 -27
rect 701 -50 703 -46
rect 748 -62 751 -39
rect 763 -54 766 -39
rect 762 -58 766 -54
rect 689 -66 691 -62
rect 747 -66 751 -62
rect 748 -71 751 -66
rect 763 -71 766 -58
rect 790 -71 792 -39
rect 865 -62 868 -39
rect 864 -66 868 -62
rect 865 -71 868 -66
rect 880 -71 883 -39
rect 907 -71 909 -39
rect 748 -81 751 -79
rect 763 -81 766 -79
rect 790 -81 792 -79
rect 865 -81 868 -79
rect 880 -81 883 -79
rect 907 -81 909 -79
rect 865 -83 872 -81
rect 869 -93 872 -83
rect 554 -97 872 -93
rect 942 -104 946 78
rect 971 74 975 165
rect 979 82 983 165
rect 1105 142 1108 146
rect 1120 142 1123 146
rect 1340 142 1343 146
rect 1355 142 1358 146
rect 1105 111 1108 134
rect 1120 119 1123 134
rect 1119 115 1123 119
rect 1104 107 1108 111
rect 1038 103 1041 107
rect 1053 103 1056 107
rect 1105 102 1108 107
rect 1120 102 1123 115
rect 1340 111 1343 134
rect 1355 119 1358 134
rect 1354 115 1358 119
rect 1173 107 1176 111
rect 1188 107 1191 111
rect 1339 107 1343 111
rect 997 86 1008 89
rect 997 -25 1000 86
rect 1005 83 1008 86
rect 1005 82 1009 83
rect 1038 72 1041 95
rect 1053 80 1056 95
rect 1273 103 1276 107
rect 1288 103 1291 107
rect 1105 92 1108 94
rect 1120 92 1123 94
rect 1052 76 1056 80
rect 1173 76 1176 99
rect 1188 84 1191 99
rect 1340 102 1343 107
rect 1355 102 1358 115
rect 1408 107 1411 111
rect 1423 107 1426 111
rect 1187 80 1191 84
rect 1037 68 1041 72
rect 1005 65 1009 66
rect 1005 23 1008 65
rect 1038 63 1041 68
rect 1053 63 1056 76
rect 1172 72 1176 76
rect 1173 67 1176 72
rect 1188 67 1191 80
rect 1105 59 1108 63
rect 1120 59 1123 63
rect 1038 53 1041 55
rect 1053 53 1056 55
rect 1173 57 1176 59
rect 1188 57 1191 59
rect 1105 28 1108 51
rect 1120 36 1123 51
rect 1119 32 1123 36
rect 1104 24 1108 28
rect 1005 20 1030 23
rect 1027 -25 1030 20
rect 1105 19 1108 24
rect 1120 19 1123 32
rect 1105 9 1108 11
rect 1120 9 1123 11
rect 997 -28 1022 -25
rect 1027 -28 1037 -25
rect 1019 -31 1022 -28
rect 1034 -31 1037 -28
rect 1061 -31 1063 -27
rect 1019 -71 1022 -39
rect 1034 -71 1037 -39
rect 1061 -71 1063 -39
rect 1019 -81 1022 -79
rect 1034 -81 1037 -79
rect 1061 -81 1063 -79
rect 1077 -93 1081 -52
rect 1212 -62 1216 -13
rect 1224 -46 1228 78
rect 1273 72 1276 95
rect 1288 80 1291 95
rect 1340 92 1343 94
rect 1355 92 1358 94
rect 1287 76 1291 80
rect 1408 76 1411 99
rect 1423 84 1426 99
rect 1422 80 1426 84
rect 1272 68 1276 72
rect 1238 -5 1242 66
rect 1273 63 1276 68
rect 1288 63 1291 76
rect 1407 72 1411 76
rect 1408 67 1411 72
rect 1423 67 1426 80
rect 1340 59 1343 63
rect 1355 59 1358 63
rect 1273 53 1276 55
rect 1288 53 1291 55
rect 1408 57 1411 59
rect 1423 57 1426 59
rect 1340 28 1343 51
rect 1355 36 1358 51
rect 1354 32 1358 36
rect 1339 24 1343 28
rect 1340 19 1343 24
rect 1355 19 1358 32
rect 1340 9 1343 11
rect 1355 9 1358 11
rect 1271 -31 1274 -27
rect 1286 -31 1289 -27
rect 1313 -31 1315 -27
rect 1388 -31 1391 -27
rect 1403 -31 1406 -27
rect 1430 -31 1432 -27
rect 1224 -50 1226 -46
rect 1271 -62 1274 -39
rect 1286 -54 1289 -39
rect 1285 -58 1289 -54
rect 1212 -66 1214 -62
rect 1270 -66 1274 -62
rect 1271 -71 1274 -66
rect 1286 -71 1289 -58
rect 1313 -71 1315 -39
rect 1388 -62 1391 -39
rect 1387 -66 1391 -62
rect 1388 -71 1391 -66
rect 1403 -71 1406 -39
rect 1430 -71 1432 -39
rect 1271 -81 1274 -79
rect 1286 -81 1289 -79
rect 1313 -81 1315 -79
rect 1388 -81 1391 -79
rect 1403 -81 1406 -79
rect 1430 -81 1432 -79
rect 1388 -83 1395 -81
rect 1392 -93 1395 -83
rect 1077 -97 1395 -93
rect 1465 -104 1469 78
<< ndiffusion >>
rect -474 100 -464 102
rect -474 96 -472 100
rect -468 96 -464 100
rect -474 94 -464 96
rect -461 94 -449 102
rect -446 100 -436 102
rect -446 96 -442 100
rect -438 96 -436 100
rect -446 94 -436 96
rect -239 100 -229 102
rect -239 96 -237 100
rect -233 96 -229 100
rect -406 65 -396 67
rect -541 61 -531 63
rect -541 57 -539 61
rect -535 57 -531 61
rect -541 55 -531 57
rect -528 55 -516 63
rect -513 61 -503 63
rect -513 57 -509 61
rect -505 57 -503 61
rect -406 61 -404 65
rect -400 61 -396 65
rect -406 59 -396 61
rect -393 59 -381 67
rect -378 65 -368 67
rect -378 61 -374 65
rect -370 61 -368 65
rect -378 59 -368 61
rect -513 55 -503 57
rect -474 17 -464 19
rect -474 13 -472 17
rect -468 13 -464 17
rect -474 11 -464 13
rect -461 11 -449 19
rect -446 17 -436 19
rect -446 13 -442 17
rect -438 13 -436 17
rect -446 11 -436 13
rect -560 -73 -550 -71
rect -560 -77 -558 -73
rect -554 -77 -550 -73
rect -560 -79 -550 -77
rect -547 -79 -535 -71
rect -532 -73 -522 -71
rect -532 -77 -528 -73
rect -524 -77 -522 -73
rect -532 -79 -522 -77
rect -518 -73 -508 -71
rect -518 -77 -516 -73
rect -512 -77 -508 -73
rect -518 -79 -508 -77
rect -506 -73 -496 -71
rect -506 -77 -502 -73
rect -498 -77 -496 -73
rect -506 -79 -496 -77
rect -239 94 -229 96
rect -226 94 -214 102
rect -211 100 -201 102
rect -211 96 -207 100
rect -203 96 -201 100
rect -211 94 -201 96
rect -171 65 -161 67
rect -306 61 -296 63
rect -306 57 -304 61
rect -300 57 -296 61
rect -306 55 -296 57
rect -293 55 -281 63
rect -278 61 -268 63
rect -278 57 -274 61
rect -270 57 -268 61
rect -171 61 -169 65
rect -165 61 -161 65
rect -171 59 -161 61
rect -158 59 -146 67
rect -143 65 -133 67
rect -143 61 -139 65
rect -135 61 -133 65
rect -143 59 -133 61
rect -278 55 -268 57
rect -239 17 -229 19
rect -239 13 -237 17
rect -233 13 -229 17
rect -239 11 -229 13
rect -226 11 -214 19
rect -211 17 -201 19
rect -211 13 -207 17
rect -203 13 -201 17
rect -211 11 -201 13
rect -308 -73 -298 -71
rect -308 -77 -306 -73
rect -302 -77 -298 -73
rect -308 -79 -298 -77
rect -295 -79 -283 -71
rect -280 -73 -270 -71
rect -280 -77 -276 -73
rect -272 -77 -270 -73
rect -280 -79 -270 -77
rect -266 -73 -256 -71
rect -266 -77 -264 -73
rect -260 -77 -256 -73
rect -266 -79 -256 -77
rect -254 -73 -244 -71
rect -254 -77 -250 -73
rect -246 -77 -244 -73
rect -254 -79 -244 -77
rect -191 -73 -181 -71
rect -191 -77 -189 -73
rect -185 -77 -181 -73
rect -191 -79 -181 -77
rect -178 -73 -166 -71
rect -178 -77 -175 -73
rect -171 -77 -166 -73
rect -178 -79 -166 -77
rect -163 -73 -153 -71
rect -163 -77 -159 -73
rect -155 -77 -153 -73
rect -163 -79 -153 -77
rect -149 -73 -139 -71
rect -149 -77 -147 -73
rect -143 -77 -139 -73
rect -149 -79 -139 -77
rect -137 -73 -127 -71
rect -137 -77 -133 -73
rect -129 -77 -127 -73
rect -137 -79 -127 -77
rect 49 100 59 102
rect 49 96 51 100
rect 55 96 59 100
rect 49 94 59 96
rect 62 94 74 102
rect 77 100 87 102
rect 77 96 81 100
rect 85 96 87 100
rect 77 94 87 96
rect 284 100 294 102
rect 284 96 286 100
rect 290 96 294 100
rect 117 65 127 67
rect -18 61 -8 63
rect -18 57 -16 61
rect -12 57 -8 61
rect -18 55 -8 57
rect -5 55 7 63
rect 10 61 20 63
rect 10 57 14 61
rect 18 57 20 61
rect 117 61 119 65
rect 123 61 127 65
rect 117 59 127 61
rect 130 59 142 67
rect 145 65 155 67
rect 145 61 149 65
rect 153 61 155 65
rect 145 59 155 61
rect 10 55 20 57
rect 49 17 59 19
rect 49 13 51 17
rect 55 13 59 17
rect 49 11 59 13
rect 62 11 74 19
rect 77 17 87 19
rect 77 13 81 17
rect 85 13 87 17
rect 77 11 87 13
rect -37 -73 -27 -71
rect -37 -77 -35 -73
rect -31 -77 -27 -73
rect -37 -79 -27 -77
rect -24 -79 -12 -71
rect -9 -73 1 -71
rect -9 -77 -5 -73
rect -1 -77 1 -73
rect -9 -79 1 -77
rect 5 -73 15 -71
rect 5 -77 7 -73
rect 11 -77 15 -73
rect 5 -79 15 -77
rect 17 -73 27 -71
rect 17 -77 21 -73
rect 25 -77 27 -73
rect 17 -79 27 -77
rect 284 94 294 96
rect 297 94 309 102
rect 312 100 322 102
rect 312 96 316 100
rect 320 96 322 100
rect 312 94 322 96
rect 352 65 362 67
rect 217 61 227 63
rect 217 57 219 61
rect 223 57 227 61
rect 217 55 227 57
rect 230 55 242 63
rect 245 61 255 63
rect 245 57 249 61
rect 253 57 255 61
rect 352 61 354 65
rect 358 61 362 65
rect 352 59 362 61
rect 365 59 377 67
rect 380 65 390 67
rect 380 61 384 65
rect 388 61 390 65
rect 380 59 390 61
rect 245 55 255 57
rect 284 17 294 19
rect 284 13 286 17
rect 290 13 294 17
rect 284 11 294 13
rect 297 11 309 19
rect 312 17 322 19
rect 312 13 316 17
rect 320 13 322 17
rect 312 11 322 13
rect 215 -73 225 -71
rect 215 -77 217 -73
rect 221 -77 225 -73
rect 215 -79 225 -77
rect 228 -79 240 -71
rect 243 -73 253 -71
rect 243 -77 247 -73
rect 251 -77 253 -73
rect 243 -79 253 -77
rect 257 -73 267 -71
rect 257 -77 259 -73
rect 263 -77 267 -73
rect 257 -79 267 -77
rect 269 -73 279 -71
rect 269 -77 273 -73
rect 277 -77 279 -73
rect 269 -79 279 -77
rect 332 -73 342 -71
rect 332 -77 334 -73
rect 338 -77 342 -73
rect 332 -79 342 -77
rect 345 -73 357 -71
rect 345 -77 348 -73
rect 352 -77 357 -73
rect 345 -79 357 -77
rect 360 -73 370 -71
rect 360 -77 364 -73
rect 368 -77 370 -73
rect 360 -79 370 -77
rect 374 -73 384 -71
rect 374 -77 376 -73
rect 380 -77 384 -73
rect 374 -79 384 -77
rect 386 -73 396 -71
rect 386 -77 390 -73
rect 394 -77 396 -73
rect 386 -79 396 -77
rect 572 100 582 102
rect 572 96 574 100
rect 578 96 582 100
rect 572 94 582 96
rect 585 94 597 102
rect 600 100 610 102
rect 600 96 604 100
rect 608 96 610 100
rect 600 94 610 96
rect 807 100 817 102
rect 807 96 809 100
rect 813 96 817 100
rect 640 65 650 67
rect 505 61 515 63
rect 505 57 507 61
rect 511 57 515 61
rect 505 55 515 57
rect 518 55 530 63
rect 533 61 543 63
rect 533 57 537 61
rect 541 57 543 61
rect 640 61 642 65
rect 646 61 650 65
rect 640 59 650 61
rect 653 59 665 67
rect 668 65 678 67
rect 668 61 672 65
rect 676 61 678 65
rect 668 59 678 61
rect 533 55 543 57
rect 572 17 582 19
rect 572 13 574 17
rect 578 13 582 17
rect 572 11 582 13
rect 585 11 597 19
rect 600 17 610 19
rect 600 13 604 17
rect 608 13 610 17
rect 600 11 610 13
rect 486 -73 496 -71
rect 486 -77 488 -73
rect 492 -77 496 -73
rect 486 -79 496 -77
rect 499 -79 511 -71
rect 514 -73 524 -71
rect 514 -77 518 -73
rect 522 -77 524 -73
rect 514 -79 524 -77
rect 528 -73 538 -71
rect 528 -77 530 -73
rect 534 -77 538 -73
rect 528 -79 538 -77
rect 540 -73 550 -71
rect 540 -77 544 -73
rect 548 -77 550 -73
rect 540 -79 550 -77
rect 807 94 817 96
rect 820 94 832 102
rect 835 100 845 102
rect 835 96 839 100
rect 843 96 845 100
rect 835 94 845 96
rect 875 65 885 67
rect 740 61 750 63
rect 740 57 742 61
rect 746 57 750 61
rect 740 55 750 57
rect 753 55 765 63
rect 768 61 778 63
rect 768 57 772 61
rect 776 57 778 61
rect 875 61 877 65
rect 881 61 885 65
rect 875 59 885 61
rect 888 59 900 67
rect 903 65 913 67
rect 903 61 907 65
rect 911 61 913 65
rect 903 59 913 61
rect 768 55 778 57
rect 807 17 817 19
rect 807 13 809 17
rect 813 13 817 17
rect 807 11 817 13
rect 820 11 832 19
rect 835 17 845 19
rect 835 13 839 17
rect 843 13 845 17
rect 835 11 845 13
rect 738 -73 748 -71
rect 738 -77 740 -73
rect 744 -77 748 -73
rect 738 -79 748 -77
rect 751 -79 763 -71
rect 766 -73 776 -71
rect 766 -77 770 -73
rect 774 -77 776 -73
rect 766 -79 776 -77
rect 780 -73 790 -71
rect 780 -77 782 -73
rect 786 -77 790 -73
rect 780 -79 790 -77
rect 792 -73 802 -71
rect 792 -77 796 -73
rect 800 -77 802 -73
rect 792 -79 802 -77
rect 855 -73 865 -71
rect 855 -77 857 -73
rect 861 -77 865 -73
rect 855 -79 865 -77
rect 868 -73 880 -71
rect 868 -77 871 -73
rect 875 -77 880 -73
rect 868 -79 880 -77
rect 883 -73 893 -71
rect 883 -77 887 -73
rect 891 -77 893 -73
rect 883 -79 893 -77
rect 897 -73 907 -71
rect 897 -77 899 -73
rect 903 -77 907 -73
rect 897 -79 907 -77
rect 909 -73 919 -71
rect 909 -77 913 -73
rect 917 -77 919 -73
rect 909 -79 919 -77
rect 1095 100 1105 102
rect 1095 96 1097 100
rect 1101 96 1105 100
rect 1095 94 1105 96
rect 1108 94 1120 102
rect 1123 100 1133 102
rect 1123 96 1127 100
rect 1131 96 1133 100
rect 1123 94 1133 96
rect 1330 100 1340 102
rect 1330 96 1332 100
rect 1336 96 1340 100
rect 1163 65 1173 67
rect 1028 61 1038 63
rect 1028 57 1030 61
rect 1034 57 1038 61
rect 1028 55 1038 57
rect 1041 55 1053 63
rect 1056 61 1066 63
rect 1056 57 1060 61
rect 1064 57 1066 61
rect 1163 61 1165 65
rect 1169 61 1173 65
rect 1163 59 1173 61
rect 1176 59 1188 67
rect 1191 65 1201 67
rect 1191 61 1195 65
rect 1199 61 1201 65
rect 1191 59 1201 61
rect 1056 55 1066 57
rect 1095 17 1105 19
rect 1095 13 1097 17
rect 1101 13 1105 17
rect 1095 11 1105 13
rect 1108 11 1120 19
rect 1123 17 1133 19
rect 1123 13 1127 17
rect 1131 13 1133 17
rect 1123 11 1133 13
rect 1009 -73 1019 -71
rect 1009 -77 1011 -73
rect 1015 -77 1019 -73
rect 1009 -79 1019 -77
rect 1022 -79 1034 -71
rect 1037 -73 1047 -71
rect 1037 -77 1041 -73
rect 1045 -77 1047 -73
rect 1037 -79 1047 -77
rect 1051 -73 1061 -71
rect 1051 -77 1053 -73
rect 1057 -77 1061 -73
rect 1051 -79 1061 -77
rect 1063 -73 1073 -71
rect 1063 -77 1067 -73
rect 1071 -77 1073 -73
rect 1063 -79 1073 -77
rect 1330 94 1340 96
rect 1343 94 1355 102
rect 1358 100 1368 102
rect 1358 96 1362 100
rect 1366 96 1368 100
rect 1358 94 1368 96
rect 1398 65 1408 67
rect 1263 61 1273 63
rect 1263 57 1265 61
rect 1269 57 1273 61
rect 1263 55 1273 57
rect 1276 55 1288 63
rect 1291 61 1301 63
rect 1291 57 1295 61
rect 1299 57 1301 61
rect 1398 61 1400 65
rect 1404 61 1408 65
rect 1398 59 1408 61
rect 1411 59 1423 67
rect 1426 65 1436 67
rect 1426 61 1430 65
rect 1434 61 1436 65
rect 1426 59 1436 61
rect 1291 55 1301 57
rect 1330 17 1340 19
rect 1330 13 1332 17
rect 1336 13 1340 17
rect 1330 11 1340 13
rect 1343 11 1355 19
rect 1358 17 1368 19
rect 1358 13 1362 17
rect 1366 13 1368 17
rect 1358 11 1368 13
rect 1261 -73 1271 -71
rect 1261 -77 1263 -73
rect 1267 -77 1271 -73
rect 1261 -79 1271 -77
rect 1274 -79 1286 -71
rect 1289 -73 1299 -71
rect 1289 -77 1293 -73
rect 1297 -77 1299 -73
rect 1289 -79 1299 -77
rect 1303 -73 1313 -71
rect 1303 -77 1305 -73
rect 1309 -77 1313 -73
rect 1303 -79 1313 -77
rect 1315 -73 1325 -71
rect 1315 -77 1319 -73
rect 1323 -77 1325 -73
rect 1315 -79 1325 -77
rect 1378 -73 1388 -71
rect 1378 -77 1380 -73
rect 1384 -77 1388 -73
rect 1378 -79 1388 -77
rect 1391 -73 1403 -71
rect 1391 -77 1394 -73
rect 1398 -77 1403 -73
rect 1391 -79 1403 -77
rect 1406 -73 1416 -71
rect 1406 -77 1410 -73
rect 1414 -77 1416 -73
rect 1406 -79 1416 -77
rect 1420 -73 1430 -71
rect 1420 -77 1422 -73
rect 1426 -77 1430 -73
rect 1420 -79 1430 -77
rect 1432 -73 1442 -71
rect 1432 -77 1436 -73
rect 1440 -77 1442 -73
rect 1432 -79 1442 -77
<< pdiffusion >>
rect -474 140 -464 142
rect -474 136 -472 140
rect -468 136 -464 140
rect -474 134 -464 136
rect -461 140 -449 142
rect -461 136 -457 140
rect -453 136 -449 140
rect -461 134 -449 136
rect -446 140 -436 142
rect -446 136 -442 140
rect -438 136 -436 140
rect -446 134 -436 136
rect -239 140 -229 142
rect -239 136 -237 140
rect -233 136 -229 140
rect -239 134 -229 136
rect -226 140 -214 142
rect -226 136 -222 140
rect -218 136 -214 140
rect -226 134 -214 136
rect -211 140 -201 142
rect -211 136 -207 140
rect -203 136 -201 140
rect -211 134 -201 136
rect -541 101 -531 103
rect -541 97 -539 101
rect -535 97 -531 101
rect -541 95 -531 97
rect -528 101 -516 103
rect -528 97 -524 101
rect -520 97 -516 101
rect -528 95 -516 97
rect -513 101 -503 103
rect -406 105 -396 107
rect -513 97 -509 101
rect -505 97 -503 101
rect -513 95 -503 97
rect -406 101 -404 105
rect -400 101 -396 105
rect -406 99 -396 101
rect -393 105 -381 107
rect -393 101 -389 105
rect -385 101 -381 105
rect -393 99 -381 101
rect -378 105 -368 107
rect -378 101 -374 105
rect -370 101 -368 105
rect -378 99 -368 101
rect -306 101 -296 103
rect -306 97 -304 101
rect -300 97 -296 101
rect -306 95 -296 97
rect -293 101 -281 103
rect -293 97 -289 101
rect -285 97 -281 101
rect -293 95 -281 97
rect -278 101 -268 103
rect -171 105 -161 107
rect -278 97 -274 101
rect -270 97 -268 101
rect -278 95 -268 97
rect -474 57 -464 59
rect -474 53 -472 57
rect -468 53 -464 57
rect -474 51 -464 53
rect -461 57 -449 59
rect -461 53 -457 57
rect -453 53 -449 57
rect -461 51 -449 53
rect -446 57 -436 59
rect -446 53 -442 57
rect -438 53 -436 57
rect -446 51 -436 53
rect -560 -33 -550 -31
rect -560 -37 -558 -33
rect -554 -37 -550 -33
rect -560 -39 -550 -37
rect -547 -33 -535 -31
rect -547 -37 -543 -33
rect -539 -37 -535 -33
rect -547 -39 -535 -37
rect -532 -33 -522 -31
rect -532 -37 -528 -33
rect -524 -37 -522 -33
rect -532 -39 -522 -37
rect -518 -33 -508 -31
rect -518 -37 -516 -33
rect -512 -37 -508 -33
rect -518 -39 -508 -37
rect -506 -33 -496 -31
rect -506 -37 -502 -33
rect -498 -37 -496 -33
rect -506 -39 -496 -37
rect -171 101 -169 105
rect -165 101 -161 105
rect -171 99 -161 101
rect -158 105 -146 107
rect -158 101 -154 105
rect -150 101 -146 105
rect -158 99 -146 101
rect -143 105 -133 107
rect -143 101 -139 105
rect -135 101 -133 105
rect -143 99 -133 101
rect -239 57 -229 59
rect -239 53 -237 57
rect -233 53 -229 57
rect -239 51 -229 53
rect -226 57 -214 59
rect -226 53 -222 57
rect -218 53 -214 57
rect -226 51 -214 53
rect -211 57 -201 59
rect -211 53 -207 57
rect -203 53 -201 57
rect -211 51 -201 53
rect -308 -33 -298 -31
rect -308 -37 -306 -33
rect -302 -37 -298 -33
rect -308 -39 -298 -37
rect -295 -33 -283 -31
rect -295 -37 -291 -33
rect -287 -37 -283 -33
rect -295 -39 -283 -37
rect -280 -33 -270 -31
rect -280 -37 -276 -33
rect -272 -37 -270 -33
rect -280 -39 -270 -37
rect -266 -33 -256 -31
rect -266 -37 -264 -33
rect -260 -37 -256 -33
rect -266 -39 -256 -37
rect -254 -33 -244 -31
rect -254 -37 -250 -33
rect -246 -37 -244 -33
rect -254 -39 -244 -37
rect -191 -33 -181 -31
rect -191 -37 -189 -33
rect -185 -37 -181 -33
rect -191 -39 -181 -37
rect -178 -39 -166 -31
rect -163 -33 -153 -31
rect -163 -37 -159 -33
rect -155 -37 -153 -33
rect -163 -39 -153 -37
rect -149 -33 -139 -31
rect -149 -37 -147 -33
rect -143 -37 -139 -33
rect -149 -39 -139 -37
rect -137 -33 -127 -31
rect -137 -37 -133 -33
rect -129 -37 -127 -33
rect -137 -39 -127 -37
rect 49 140 59 142
rect 49 136 51 140
rect 55 136 59 140
rect 49 134 59 136
rect 62 140 74 142
rect 62 136 66 140
rect 70 136 74 140
rect 62 134 74 136
rect 77 140 87 142
rect 77 136 81 140
rect 85 136 87 140
rect 77 134 87 136
rect 284 140 294 142
rect 284 136 286 140
rect 290 136 294 140
rect 284 134 294 136
rect 297 140 309 142
rect 297 136 301 140
rect 305 136 309 140
rect 297 134 309 136
rect 312 140 322 142
rect 312 136 316 140
rect 320 136 322 140
rect 312 134 322 136
rect -18 101 -8 103
rect -18 97 -16 101
rect -12 97 -8 101
rect -18 95 -8 97
rect -5 101 7 103
rect -5 97 -1 101
rect 3 97 7 101
rect -5 95 7 97
rect 10 101 20 103
rect 117 105 127 107
rect 10 97 14 101
rect 18 97 20 101
rect 10 95 20 97
rect 117 101 119 105
rect 123 101 127 105
rect 117 99 127 101
rect 130 105 142 107
rect 130 101 134 105
rect 138 101 142 105
rect 130 99 142 101
rect 145 105 155 107
rect 145 101 149 105
rect 153 101 155 105
rect 145 99 155 101
rect 217 101 227 103
rect 217 97 219 101
rect 223 97 227 101
rect 217 95 227 97
rect 230 101 242 103
rect 230 97 234 101
rect 238 97 242 101
rect 230 95 242 97
rect 245 101 255 103
rect 352 105 362 107
rect 245 97 249 101
rect 253 97 255 101
rect 245 95 255 97
rect 49 57 59 59
rect 49 53 51 57
rect 55 53 59 57
rect 49 51 59 53
rect 62 57 74 59
rect 62 53 66 57
rect 70 53 74 57
rect 62 51 74 53
rect 77 57 87 59
rect 77 53 81 57
rect 85 53 87 57
rect 77 51 87 53
rect -37 -33 -27 -31
rect -37 -37 -35 -33
rect -31 -37 -27 -33
rect -37 -39 -27 -37
rect -24 -33 -12 -31
rect -24 -37 -20 -33
rect -16 -37 -12 -33
rect -24 -39 -12 -37
rect -9 -33 1 -31
rect -9 -37 -5 -33
rect -1 -37 1 -33
rect -9 -39 1 -37
rect 5 -33 15 -31
rect 5 -37 7 -33
rect 11 -37 15 -33
rect 5 -39 15 -37
rect 17 -33 27 -31
rect 17 -37 21 -33
rect 25 -37 27 -33
rect 17 -39 27 -37
rect 352 101 354 105
rect 358 101 362 105
rect 352 99 362 101
rect 365 105 377 107
rect 365 101 369 105
rect 373 101 377 105
rect 365 99 377 101
rect 380 105 390 107
rect 380 101 384 105
rect 388 101 390 105
rect 380 99 390 101
rect 284 57 294 59
rect 284 53 286 57
rect 290 53 294 57
rect 284 51 294 53
rect 297 57 309 59
rect 297 53 301 57
rect 305 53 309 57
rect 297 51 309 53
rect 312 57 322 59
rect 312 53 316 57
rect 320 53 322 57
rect 312 51 322 53
rect 215 -33 225 -31
rect 215 -37 217 -33
rect 221 -37 225 -33
rect 215 -39 225 -37
rect 228 -33 240 -31
rect 228 -37 232 -33
rect 236 -37 240 -33
rect 228 -39 240 -37
rect 243 -33 253 -31
rect 243 -37 247 -33
rect 251 -37 253 -33
rect 243 -39 253 -37
rect 257 -33 267 -31
rect 257 -37 259 -33
rect 263 -37 267 -33
rect 257 -39 267 -37
rect 269 -33 279 -31
rect 269 -37 273 -33
rect 277 -37 279 -33
rect 269 -39 279 -37
rect 332 -33 342 -31
rect 332 -37 334 -33
rect 338 -37 342 -33
rect 332 -39 342 -37
rect 345 -39 357 -31
rect 360 -33 370 -31
rect 360 -37 364 -33
rect 368 -37 370 -33
rect 360 -39 370 -37
rect 374 -33 384 -31
rect 374 -37 376 -33
rect 380 -37 384 -33
rect 374 -39 384 -37
rect 386 -33 396 -31
rect 386 -37 390 -33
rect 394 -37 396 -33
rect 386 -39 396 -37
rect 572 140 582 142
rect 572 136 574 140
rect 578 136 582 140
rect 572 134 582 136
rect 585 140 597 142
rect 585 136 589 140
rect 593 136 597 140
rect 585 134 597 136
rect 600 140 610 142
rect 600 136 604 140
rect 608 136 610 140
rect 600 134 610 136
rect 807 140 817 142
rect 807 136 809 140
rect 813 136 817 140
rect 807 134 817 136
rect 820 140 832 142
rect 820 136 824 140
rect 828 136 832 140
rect 820 134 832 136
rect 835 140 845 142
rect 835 136 839 140
rect 843 136 845 140
rect 835 134 845 136
rect 505 101 515 103
rect 505 97 507 101
rect 511 97 515 101
rect 505 95 515 97
rect 518 101 530 103
rect 518 97 522 101
rect 526 97 530 101
rect 518 95 530 97
rect 533 101 543 103
rect 640 105 650 107
rect 533 97 537 101
rect 541 97 543 101
rect 533 95 543 97
rect 640 101 642 105
rect 646 101 650 105
rect 640 99 650 101
rect 653 105 665 107
rect 653 101 657 105
rect 661 101 665 105
rect 653 99 665 101
rect 668 105 678 107
rect 668 101 672 105
rect 676 101 678 105
rect 668 99 678 101
rect 740 101 750 103
rect 740 97 742 101
rect 746 97 750 101
rect 740 95 750 97
rect 753 101 765 103
rect 753 97 757 101
rect 761 97 765 101
rect 753 95 765 97
rect 768 101 778 103
rect 875 105 885 107
rect 768 97 772 101
rect 776 97 778 101
rect 768 95 778 97
rect 572 57 582 59
rect 572 53 574 57
rect 578 53 582 57
rect 572 51 582 53
rect 585 57 597 59
rect 585 53 589 57
rect 593 53 597 57
rect 585 51 597 53
rect 600 57 610 59
rect 600 53 604 57
rect 608 53 610 57
rect 600 51 610 53
rect 486 -33 496 -31
rect 486 -37 488 -33
rect 492 -37 496 -33
rect 486 -39 496 -37
rect 499 -33 511 -31
rect 499 -37 503 -33
rect 507 -37 511 -33
rect 499 -39 511 -37
rect 514 -33 524 -31
rect 514 -37 518 -33
rect 522 -37 524 -33
rect 514 -39 524 -37
rect 528 -33 538 -31
rect 528 -37 530 -33
rect 534 -37 538 -33
rect 528 -39 538 -37
rect 540 -33 550 -31
rect 540 -37 544 -33
rect 548 -37 550 -33
rect 540 -39 550 -37
rect 875 101 877 105
rect 881 101 885 105
rect 875 99 885 101
rect 888 105 900 107
rect 888 101 892 105
rect 896 101 900 105
rect 888 99 900 101
rect 903 105 913 107
rect 903 101 907 105
rect 911 101 913 105
rect 903 99 913 101
rect 807 57 817 59
rect 807 53 809 57
rect 813 53 817 57
rect 807 51 817 53
rect 820 57 832 59
rect 820 53 824 57
rect 828 53 832 57
rect 820 51 832 53
rect 835 57 845 59
rect 835 53 839 57
rect 843 53 845 57
rect 835 51 845 53
rect 738 -33 748 -31
rect 738 -37 740 -33
rect 744 -37 748 -33
rect 738 -39 748 -37
rect 751 -33 763 -31
rect 751 -37 755 -33
rect 759 -37 763 -33
rect 751 -39 763 -37
rect 766 -33 776 -31
rect 766 -37 770 -33
rect 774 -37 776 -33
rect 766 -39 776 -37
rect 780 -33 790 -31
rect 780 -37 782 -33
rect 786 -37 790 -33
rect 780 -39 790 -37
rect 792 -33 802 -31
rect 792 -37 796 -33
rect 800 -37 802 -33
rect 792 -39 802 -37
rect 855 -33 865 -31
rect 855 -37 857 -33
rect 861 -37 865 -33
rect 855 -39 865 -37
rect 868 -39 880 -31
rect 883 -33 893 -31
rect 883 -37 887 -33
rect 891 -37 893 -33
rect 883 -39 893 -37
rect 897 -33 907 -31
rect 897 -37 899 -33
rect 903 -37 907 -33
rect 897 -39 907 -37
rect 909 -33 919 -31
rect 909 -37 913 -33
rect 917 -37 919 -33
rect 909 -39 919 -37
rect 1095 140 1105 142
rect 1095 136 1097 140
rect 1101 136 1105 140
rect 1095 134 1105 136
rect 1108 140 1120 142
rect 1108 136 1112 140
rect 1116 136 1120 140
rect 1108 134 1120 136
rect 1123 140 1133 142
rect 1123 136 1127 140
rect 1131 136 1133 140
rect 1123 134 1133 136
rect 1330 140 1340 142
rect 1330 136 1332 140
rect 1336 136 1340 140
rect 1330 134 1340 136
rect 1343 140 1355 142
rect 1343 136 1347 140
rect 1351 136 1355 140
rect 1343 134 1355 136
rect 1358 140 1368 142
rect 1358 136 1362 140
rect 1366 136 1368 140
rect 1358 134 1368 136
rect 1028 101 1038 103
rect 1028 97 1030 101
rect 1034 97 1038 101
rect 1028 95 1038 97
rect 1041 101 1053 103
rect 1041 97 1045 101
rect 1049 97 1053 101
rect 1041 95 1053 97
rect 1056 101 1066 103
rect 1163 105 1173 107
rect 1056 97 1060 101
rect 1064 97 1066 101
rect 1056 95 1066 97
rect 1163 101 1165 105
rect 1169 101 1173 105
rect 1163 99 1173 101
rect 1176 105 1188 107
rect 1176 101 1180 105
rect 1184 101 1188 105
rect 1176 99 1188 101
rect 1191 105 1201 107
rect 1191 101 1195 105
rect 1199 101 1201 105
rect 1191 99 1201 101
rect 1263 101 1273 103
rect 1263 97 1265 101
rect 1269 97 1273 101
rect 1263 95 1273 97
rect 1276 101 1288 103
rect 1276 97 1280 101
rect 1284 97 1288 101
rect 1276 95 1288 97
rect 1291 101 1301 103
rect 1398 105 1408 107
rect 1291 97 1295 101
rect 1299 97 1301 101
rect 1291 95 1301 97
rect 1095 57 1105 59
rect 1095 53 1097 57
rect 1101 53 1105 57
rect 1095 51 1105 53
rect 1108 57 1120 59
rect 1108 53 1112 57
rect 1116 53 1120 57
rect 1108 51 1120 53
rect 1123 57 1133 59
rect 1123 53 1127 57
rect 1131 53 1133 57
rect 1123 51 1133 53
rect 1009 -33 1019 -31
rect 1009 -37 1011 -33
rect 1015 -37 1019 -33
rect 1009 -39 1019 -37
rect 1022 -33 1034 -31
rect 1022 -37 1026 -33
rect 1030 -37 1034 -33
rect 1022 -39 1034 -37
rect 1037 -33 1047 -31
rect 1037 -37 1041 -33
rect 1045 -37 1047 -33
rect 1037 -39 1047 -37
rect 1051 -33 1061 -31
rect 1051 -37 1053 -33
rect 1057 -37 1061 -33
rect 1051 -39 1061 -37
rect 1063 -33 1073 -31
rect 1063 -37 1067 -33
rect 1071 -37 1073 -33
rect 1063 -39 1073 -37
rect 1398 101 1400 105
rect 1404 101 1408 105
rect 1398 99 1408 101
rect 1411 105 1423 107
rect 1411 101 1415 105
rect 1419 101 1423 105
rect 1411 99 1423 101
rect 1426 105 1436 107
rect 1426 101 1430 105
rect 1434 101 1436 105
rect 1426 99 1436 101
rect 1330 57 1340 59
rect 1330 53 1332 57
rect 1336 53 1340 57
rect 1330 51 1340 53
rect 1343 57 1355 59
rect 1343 53 1347 57
rect 1351 53 1355 57
rect 1343 51 1355 53
rect 1358 57 1368 59
rect 1358 53 1362 57
rect 1366 53 1368 57
rect 1358 51 1368 53
rect 1261 -33 1271 -31
rect 1261 -37 1263 -33
rect 1267 -37 1271 -33
rect 1261 -39 1271 -37
rect 1274 -33 1286 -31
rect 1274 -37 1278 -33
rect 1282 -37 1286 -33
rect 1274 -39 1286 -37
rect 1289 -33 1299 -31
rect 1289 -37 1293 -33
rect 1297 -37 1299 -33
rect 1289 -39 1299 -37
rect 1303 -33 1313 -31
rect 1303 -37 1305 -33
rect 1309 -37 1313 -33
rect 1303 -39 1313 -37
rect 1315 -33 1325 -31
rect 1315 -37 1319 -33
rect 1323 -37 1325 -33
rect 1315 -39 1325 -37
rect 1378 -33 1388 -31
rect 1378 -37 1380 -33
rect 1384 -37 1388 -33
rect 1378 -39 1388 -37
rect 1391 -39 1403 -31
rect 1406 -33 1416 -31
rect 1406 -37 1410 -33
rect 1414 -37 1416 -33
rect 1406 -39 1416 -37
rect 1420 -33 1430 -31
rect 1420 -37 1422 -33
rect 1426 -37 1430 -33
rect 1420 -39 1430 -37
rect 1432 -33 1442 -31
rect 1432 -37 1436 -33
rect 1440 -37 1442 -33
rect 1432 -39 1442 -37
<< metal1 >>
rect -612 152 -467 154
rect -612 150 -504 152
rect -500 150 -467 152
rect -463 150 -448 154
rect -444 152 -232 154
rect -444 150 -269 152
rect -472 140 -468 150
rect -442 140 -438 150
rect -457 127 -453 136
rect -457 123 -438 127
rect -551 119 -476 123
rect -442 119 -438 123
rect -387 119 -383 150
rect -265 150 -232 152
rect -228 150 -213 154
rect -209 152 56 154
rect -209 150 -113 152
rect -237 140 -233 150
rect -207 140 -203 150
rect -222 127 -218 136
rect -222 123 -203 127
rect -316 119 -241 123
rect -207 119 -203 123
rect -152 119 -148 150
rect -109 150 19 152
rect 23 150 56 152
rect 60 150 75 154
rect 79 152 291 154
rect 79 150 254 152
rect 51 140 55 150
rect 81 140 85 150
rect 66 127 70 136
rect 66 123 85 127
rect -28 119 47 123
rect 81 119 85 123
rect 136 119 140 150
rect 258 150 291 152
rect 295 150 310 154
rect 314 152 579 154
rect 314 150 410 152
rect 286 140 290 150
rect 316 140 320 150
rect 301 127 305 136
rect 301 123 320 127
rect 207 119 282 123
rect 316 119 320 123
rect 371 119 375 150
rect 414 150 542 152
rect 546 150 579 152
rect 583 150 598 154
rect 602 152 814 154
rect 602 150 777 152
rect 574 140 578 150
rect 604 140 608 150
rect 589 127 593 136
rect 589 123 608 127
rect 495 119 570 123
rect 604 119 608 123
rect 659 119 663 150
rect 781 150 814 152
rect 818 150 833 154
rect 837 152 1102 154
rect 837 150 933 152
rect 809 140 813 150
rect 839 140 843 150
rect 824 127 828 136
rect 824 123 843 127
rect 730 119 805 123
rect 839 119 843 123
rect 894 119 898 150
rect 937 150 1065 152
rect 1069 150 1102 152
rect 1106 150 1121 154
rect 1125 152 1337 154
rect 1125 150 1300 152
rect 1097 140 1101 150
rect 1127 140 1131 150
rect 1112 127 1116 136
rect 1112 123 1131 127
rect 1018 119 1093 123
rect 1127 119 1131 123
rect 1182 119 1186 150
rect 1304 150 1337 152
rect 1341 150 1356 154
rect 1360 152 1480 154
rect 1360 150 1456 152
rect 1332 140 1336 150
rect 1362 140 1366 150
rect 1347 127 1351 136
rect 1347 123 1366 127
rect 1253 119 1328 123
rect 1362 119 1366 123
rect 1417 119 1421 150
rect 1460 150 1480 152
rect -586 78 -564 80
rect -551 80 -546 119
rect -480 115 -454 119
rect -442 115 -422 119
rect -406 115 -399 119
rect -395 115 -380 119
rect -376 115 -366 119
rect -543 111 -534 115
rect -530 111 -515 115
rect -511 111 -506 115
rect -539 101 -535 111
rect -509 101 -505 111
rect -489 107 -469 111
rect -524 88 -520 97
rect -524 84 -505 88
rect -509 80 -505 84
rect -489 80 -485 107
rect -442 100 -438 115
rect -472 88 -468 96
rect -474 84 -467 88
rect -463 84 -446 88
rect -442 84 -438 88
rect -426 84 -422 115
rect -404 105 -400 115
rect -374 105 -370 115
rect -389 92 -385 101
rect -389 88 -370 92
rect -374 84 -370 88
rect -316 84 -311 119
rect -245 115 -219 119
rect -207 115 -187 119
rect -171 115 -164 119
rect -160 115 -145 119
rect -141 115 -131 119
rect -308 111 -299 115
rect -295 111 -280 115
rect -276 111 -271 115
rect -304 101 -300 111
rect -274 101 -270 111
rect -254 107 -234 111
rect -289 88 -285 97
rect -289 84 -270 88
rect -426 80 -386 84
rect -374 82 -311 84
rect -374 80 -345 82
rect -560 78 -521 80
rect -590 76 -521 78
rect -509 76 -485 80
rect -600 70 -598 72
rect -594 70 -536 72
rect -600 68 -564 70
rect -560 68 -536 70
rect -549 41 -544 68
rect -509 61 -505 76
rect -539 49 -535 57
rect -541 45 -534 49
rect -530 45 -513 49
rect -509 45 -504 49
rect -549 37 -494 41
rect -499 28 -494 37
rect -489 36 -485 76
rect -426 72 -401 76
rect -473 67 -467 71
rect -463 67 -448 71
rect -444 67 -436 71
rect -472 57 -468 67
rect -442 57 -438 67
rect -457 44 -453 53
rect -457 40 -438 44
rect -442 36 -438 40
rect -426 36 -422 72
rect -374 65 -370 80
rect -341 80 -311 82
rect -274 80 -270 84
rect -254 80 -250 107
rect -207 100 -203 115
rect -237 88 -233 96
rect -239 84 -232 88
rect -228 84 -211 88
rect -207 84 -203 88
rect -191 84 -187 115
rect -169 105 -165 115
rect -139 105 -135 115
rect -154 92 -150 101
rect -154 88 -135 92
rect -139 84 -135 88
rect -191 80 -151 84
rect -139 82 -100 84
rect -139 80 -104 82
rect -316 76 -286 80
rect -274 76 -250 80
rect -331 70 -301 72
rect -327 68 -301 70
rect -404 53 -400 61
rect -404 49 -399 53
rect -395 49 -378 53
rect -374 49 -370 53
rect -314 41 -309 68
rect -274 61 -270 76
rect -304 49 -300 57
rect -306 45 -299 49
rect -295 45 -278 49
rect -274 45 -269 49
rect -314 37 -259 41
rect -489 32 -454 36
rect -442 32 -422 36
rect -499 24 -469 28
rect -442 17 -438 32
rect -264 28 -259 37
rect -254 36 -250 76
rect -191 72 -166 76
rect -238 67 -232 71
rect -228 67 -213 71
rect -209 67 -201 71
rect -237 57 -233 67
rect -207 57 -203 67
rect -222 44 -218 53
rect -222 40 -203 44
rect -207 36 -203 40
rect -191 36 -187 72
rect -139 65 -135 80
rect -63 78 -41 80
rect -28 80 -23 119
rect 43 115 69 119
rect 81 115 101 119
rect 117 115 124 119
rect 128 115 143 119
rect 147 115 157 119
rect -20 111 -11 115
rect -7 111 8 115
rect 12 111 17 115
rect -16 101 -12 111
rect 14 101 18 111
rect 34 107 54 111
rect -1 88 3 97
rect -1 84 18 88
rect 14 80 18 84
rect 34 80 38 107
rect 81 100 85 115
rect 51 88 55 96
rect 49 84 56 88
rect 60 84 77 88
rect 81 84 85 88
rect 97 84 101 115
rect 119 105 123 115
rect 149 105 153 115
rect 134 92 138 101
rect 134 88 153 92
rect 149 84 153 88
rect 207 84 212 119
rect 278 115 304 119
rect 316 115 336 119
rect 352 115 359 119
rect 363 115 378 119
rect 382 115 392 119
rect 215 111 224 115
rect 228 111 243 115
rect 247 111 252 115
rect 219 101 223 111
rect 249 101 253 111
rect 269 107 289 111
rect 234 88 238 97
rect 234 84 253 88
rect 97 80 137 84
rect 149 82 212 84
rect 149 80 178 82
rect -37 78 2 80
rect -67 76 2 78
rect 14 76 38 80
rect -77 70 -75 72
rect -71 70 -13 72
rect -77 68 -41 70
rect -37 68 -13 70
rect -169 53 -165 61
rect -169 49 -164 53
rect -160 49 -143 53
rect -139 49 -135 53
rect -26 41 -21 68
rect 14 61 18 76
rect -16 49 -12 57
rect -18 45 -11 49
rect -7 45 10 49
rect 14 45 19 49
rect -26 37 29 41
rect -254 32 -219 36
rect -207 32 -187 36
rect -264 24 -234 28
rect -207 17 -203 32
rect 24 28 29 37
rect 34 36 38 76
rect 97 72 122 76
rect 50 67 56 71
rect 60 67 75 71
rect 79 67 87 71
rect 51 57 55 67
rect 81 57 85 67
rect 66 44 70 53
rect 66 40 85 44
rect 81 36 85 40
rect 97 36 101 72
rect 149 65 153 80
rect 182 80 212 82
rect 249 80 253 84
rect 269 80 273 107
rect 316 100 320 115
rect 286 88 290 96
rect 284 84 291 88
rect 295 84 312 88
rect 316 84 320 88
rect 332 84 336 115
rect 354 105 358 115
rect 384 105 388 115
rect 369 92 373 101
rect 369 88 388 92
rect 384 84 388 88
rect 332 80 372 84
rect 384 82 423 84
rect 384 80 419 82
rect 207 76 237 80
rect 249 76 273 80
rect 192 70 222 72
rect 196 68 222 70
rect 119 53 123 61
rect 119 49 124 53
rect 128 49 145 53
rect 149 49 153 53
rect 209 41 214 68
rect 249 61 253 76
rect 219 49 223 57
rect 217 45 224 49
rect 228 45 245 49
rect 249 45 254 49
rect 209 37 264 41
rect 34 32 69 36
rect 81 32 101 36
rect 24 24 54 28
rect 81 17 85 32
rect 259 28 264 37
rect 269 36 273 76
rect 332 72 357 76
rect 285 67 291 71
rect 295 67 310 71
rect 314 67 322 71
rect 286 57 290 67
rect 316 57 320 67
rect 301 44 305 53
rect 301 40 320 44
rect 316 36 320 40
rect 332 36 336 72
rect 384 65 388 80
rect 460 78 482 80
rect 495 80 500 119
rect 566 115 592 119
rect 604 115 624 119
rect 640 115 647 119
rect 651 115 666 119
rect 670 115 680 119
rect 503 111 512 115
rect 516 111 531 115
rect 535 111 540 115
rect 507 101 511 111
rect 537 101 541 111
rect 557 107 577 111
rect 522 88 526 97
rect 522 84 541 88
rect 537 80 541 84
rect 557 80 561 107
rect 604 100 608 115
rect 574 88 578 96
rect 572 84 579 88
rect 583 84 600 88
rect 604 84 608 88
rect 620 84 624 115
rect 642 105 646 115
rect 672 105 676 115
rect 657 92 661 101
rect 657 88 676 92
rect 672 84 676 88
rect 730 84 735 119
rect 801 115 827 119
rect 839 115 859 119
rect 875 115 882 119
rect 886 115 901 119
rect 905 115 915 119
rect 738 111 747 115
rect 751 111 766 115
rect 770 111 775 115
rect 742 101 746 111
rect 772 101 776 111
rect 792 107 812 111
rect 757 88 761 97
rect 757 84 776 88
rect 620 80 660 84
rect 672 82 735 84
rect 672 80 701 82
rect 486 78 525 80
rect 456 76 525 78
rect 537 76 561 80
rect 446 70 448 72
rect 452 70 510 72
rect 446 68 482 70
rect 486 68 510 70
rect 354 53 358 61
rect 354 49 359 53
rect 363 49 380 53
rect 384 49 388 53
rect 497 41 502 68
rect 537 61 541 76
rect 507 49 511 57
rect 505 45 512 49
rect 516 45 533 49
rect 537 45 542 49
rect 497 37 552 41
rect 269 32 304 36
rect 316 32 336 36
rect 259 24 289 28
rect 316 17 320 32
rect 547 28 552 37
rect 557 36 561 76
rect 620 72 645 76
rect 573 67 579 71
rect 583 67 598 71
rect 602 67 610 71
rect 574 57 578 67
rect 604 57 608 67
rect 589 44 593 53
rect 589 40 608 44
rect 604 36 608 40
rect 620 36 624 72
rect 672 65 676 80
rect 705 80 735 82
rect 772 80 776 84
rect 792 80 796 107
rect 839 100 843 115
rect 809 88 813 96
rect 807 84 814 88
rect 818 84 835 88
rect 839 84 843 88
rect 855 84 859 115
rect 877 105 881 115
rect 907 105 911 115
rect 892 92 896 101
rect 892 88 911 92
rect 907 84 911 88
rect 855 80 895 84
rect 907 82 946 84
rect 907 80 942 82
rect 730 76 760 80
rect 772 76 796 80
rect 715 70 745 72
rect 719 68 745 70
rect 642 53 646 61
rect 642 49 647 53
rect 651 49 668 53
rect 672 49 676 53
rect 732 41 737 68
rect 772 61 776 76
rect 742 49 746 57
rect 740 45 747 49
rect 751 45 768 49
rect 772 45 777 49
rect 732 37 787 41
rect 557 32 592 36
rect 604 32 624 36
rect 547 24 577 28
rect 604 17 608 32
rect 782 28 787 37
rect 792 36 796 76
rect 855 72 880 76
rect 808 67 814 71
rect 818 67 833 71
rect 837 67 845 71
rect 809 57 813 67
rect 839 57 843 67
rect 824 44 828 53
rect 824 40 843 44
rect 839 36 843 40
rect 855 36 859 72
rect 907 65 911 80
rect 983 78 1005 80
rect 1018 80 1023 119
rect 1089 115 1115 119
rect 1127 115 1147 119
rect 1163 115 1170 119
rect 1174 115 1189 119
rect 1193 115 1203 119
rect 1026 111 1035 115
rect 1039 111 1054 115
rect 1058 111 1063 115
rect 1030 101 1034 111
rect 1060 101 1064 111
rect 1080 107 1100 111
rect 1045 88 1049 97
rect 1045 84 1064 88
rect 1060 80 1064 84
rect 1080 80 1084 107
rect 1127 100 1131 115
rect 1097 88 1101 96
rect 1095 84 1102 88
rect 1106 84 1123 88
rect 1127 84 1131 88
rect 1143 84 1147 115
rect 1165 105 1169 115
rect 1195 105 1199 115
rect 1180 92 1184 101
rect 1180 88 1199 92
rect 1195 84 1199 88
rect 1253 84 1258 119
rect 1324 115 1350 119
rect 1362 115 1382 119
rect 1398 115 1405 119
rect 1409 115 1424 119
rect 1428 115 1438 119
rect 1261 111 1270 115
rect 1274 111 1289 115
rect 1293 111 1298 115
rect 1265 101 1269 111
rect 1295 101 1299 111
rect 1315 107 1335 111
rect 1280 88 1284 97
rect 1280 84 1299 88
rect 1143 80 1183 84
rect 1195 82 1258 84
rect 1195 80 1224 82
rect 1009 78 1048 80
rect 979 76 1048 78
rect 1060 76 1084 80
rect 969 70 971 72
rect 975 70 1033 72
rect 969 68 1005 70
rect 1009 68 1033 70
rect 877 53 881 61
rect 877 49 882 53
rect 886 49 903 53
rect 907 49 911 53
rect 1020 41 1025 68
rect 1060 61 1064 76
rect 1030 49 1034 57
rect 1028 45 1035 49
rect 1039 45 1056 49
rect 1060 45 1065 49
rect 1020 37 1075 41
rect 792 32 827 36
rect 839 32 859 36
rect 782 24 812 28
rect 839 17 843 32
rect 1070 28 1075 37
rect 1080 36 1084 76
rect 1143 72 1168 76
rect 1096 67 1102 71
rect 1106 67 1121 71
rect 1125 67 1133 71
rect 1097 57 1101 67
rect 1127 57 1131 67
rect 1112 44 1116 53
rect 1112 40 1131 44
rect 1127 36 1131 40
rect 1143 36 1147 72
rect 1195 65 1199 80
rect 1228 80 1258 82
rect 1295 80 1299 84
rect 1315 80 1319 107
rect 1362 100 1366 115
rect 1332 88 1336 96
rect 1330 84 1337 88
rect 1341 84 1358 88
rect 1362 84 1366 88
rect 1378 84 1382 115
rect 1400 105 1404 115
rect 1430 105 1434 115
rect 1415 92 1419 101
rect 1415 88 1434 92
rect 1430 84 1434 88
rect 1378 80 1418 84
rect 1430 82 1469 84
rect 1430 80 1465 82
rect 1253 76 1283 80
rect 1295 76 1319 80
rect 1238 70 1268 72
rect 1242 68 1268 70
rect 1165 53 1169 61
rect 1165 49 1170 53
rect 1174 49 1191 53
rect 1195 49 1199 53
rect 1255 41 1260 68
rect 1295 61 1299 76
rect 1265 49 1269 57
rect 1263 45 1270 49
rect 1274 45 1291 49
rect 1295 45 1300 49
rect 1255 37 1310 41
rect 1080 32 1115 36
rect 1127 32 1147 36
rect 1070 24 1100 28
rect 1127 17 1131 32
rect 1305 28 1310 37
rect 1315 36 1319 76
rect 1378 72 1403 76
rect 1331 67 1337 71
rect 1341 67 1356 71
rect 1360 67 1368 71
rect 1332 57 1336 67
rect 1362 57 1366 67
rect 1347 44 1351 53
rect 1347 40 1366 44
rect 1362 36 1366 40
rect 1378 36 1382 72
rect 1430 65 1434 80
rect 1400 53 1404 61
rect 1400 49 1405 53
rect 1409 49 1426 53
rect 1430 49 1434 53
rect 1315 32 1350 36
rect 1362 32 1382 36
rect 1305 24 1335 28
rect 1362 17 1366 32
rect -505 3 -494 5
rect -472 5 -468 13
rect -490 3 -467 5
rect -505 1 -467 3
rect -463 1 -446 5
rect -442 3 -434 5
rect -430 3 -410 5
rect -406 3 -259 5
rect -237 5 -233 13
rect -255 3 -232 5
rect -442 1 -232 3
rect -228 1 -211 5
rect -207 3 -199 5
rect -195 3 -175 5
rect -171 3 -107 5
rect -207 1 -121 3
rect -117 1 -107 3
rect 18 3 29 5
rect 51 5 55 13
rect 33 3 56 5
rect 18 1 56 3
rect 60 1 77 5
rect 81 3 89 5
rect 93 3 113 5
rect 117 3 264 5
rect 286 5 290 13
rect 268 3 291 5
rect 81 1 291 3
rect 295 1 312 5
rect 316 3 324 5
rect 328 3 348 5
rect 352 3 416 5
rect 316 1 402 3
rect 406 1 416 3
rect 541 3 552 5
rect 574 5 578 13
rect 556 3 579 5
rect 541 1 579 3
rect 583 1 600 5
rect 604 3 612 5
rect 616 3 636 5
rect 640 3 787 5
rect 809 5 813 13
rect 791 3 814 5
rect 604 1 814 3
rect 818 1 835 5
rect 839 3 847 5
rect 851 3 871 5
rect 875 3 939 5
rect 839 1 925 3
rect 929 1 939 3
rect 1064 3 1075 5
rect 1097 5 1101 13
rect 1079 3 1102 5
rect 1064 1 1102 3
rect 1106 1 1123 5
rect 1127 3 1135 5
rect 1139 3 1159 5
rect 1163 3 1310 5
rect 1332 5 1336 13
rect 1314 3 1337 5
rect 1127 1 1337 3
rect 1341 1 1358 5
rect 1362 3 1370 5
rect 1374 3 1394 5
rect 1398 3 1462 5
rect 1362 1 1448 3
rect 1452 1 1462 3
rect -601 -9 -331 -7
rect -601 -11 -357 -9
rect -601 -52 -597 -11
rect -353 -11 -327 -9
rect -78 -9 192 -7
rect -78 -11 166 -9
rect -561 -23 -553 -19
rect -549 -23 -534 -19
rect -530 -23 -516 -19
rect -512 -23 -502 -19
rect -498 -23 -301 -19
rect -297 -23 -282 -19
rect -278 -23 -264 -19
rect -260 -23 -250 -19
rect -246 -23 -184 -19
rect -180 -23 -165 -19
rect -161 -23 -147 -19
rect -143 -23 -133 -19
rect -129 -21 -113 -19
rect -109 -21 -107 -19
rect -129 -23 -107 -21
rect -558 -33 -554 -23
rect -528 -33 -524 -23
rect -516 -33 -512 -23
rect -306 -33 -302 -23
rect -276 -33 -272 -23
rect -264 -33 -260 -23
rect -189 -33 -185 -23
rect -147 -33 -143 -23
rect -543 -46 -539 -37
rect -543 -50 -524 -46
rect -612 -56 -597 -52
rect -528 -54 -524 -50
rect -502 -52 -498 -37
rect -291 -46 -287 -37
rect -250 -46 -246 -37
rect -339 -50 -299 -46
rect -291 -50 -272 -46
rect -528 -58 -512 -54
rect -502 -56 -496 -52
rect -303 -54 -299 -50
rect -276 -54 -272 -50
rect -250 -50 -170 -46
rect -528 -73 -524 -58
rect -502 -73 -498 -56
rect -303 -58 -288 -54
rect -276 -58 -260 -54
rect -351 -66 -303 -62
rect -276 -73 -272 -58
rect -250 -73 -246 -50
rect -159 -54 -155 -37
rect -133 -52 -129 -37
rect -78 -52 -74 -11
rect 170 -11 196 -9
rect 445 -9 715 -7
rect 445 -11 689 -9
rect -38 -23 -30 -19
rect -26 -23 -11 -19
rect -7 -23 7 -19
rect 11 -23 21 -19
rect 25 -23 222 -19
rect 226 -23 241 -19
rect 245 -23 259 -19
rect 263 -23 273 -19
rect 277 -23 339 -19
rect 343 -23 358 -19
rect 362 -23 376 -19
rect 380 -23 390 -19
rect 394 -21 410 -19
rect 414 -21 416 -19
rect 394 -23 416 -21
rect -35 -33 -31 -23
rect -5 -33 -1 -23
rect 7 -33 11 -23
rect 217 -33 221 -23
rect 247 -33 251 -23
rect 259 -33 263 -23
rect 334 -33 338 -23
rect 376 -33 380 -23
rect -20 -46 -16 -37
rect -20 -50 -1 -46
rect -175 -58 -143 -54
rect -133 -56 -74 -52
rect -5 -54 -1 -50
rect 21 -52 25 -37
rect 232 -46 236 -37
rect 273 -46 277 -37
rect 184 -50 224 -46
rect 232 -50 251 -46
rect -193 -66 -186 -62
rect -175 -73 -171 -58
rect -133 -73 -129 -56
rect -5 -58 11 -54
rect 21 -56 27 -52
rect 220 -54 224 -50
rect 247 -54 251 -50
rect 273 -50 353 -46
rect -5 -73 -1 -58
rect 21 -73 25 -56
rect 220 -58 235 -54
rect 247 -58 263 -54
rect 172 -66 220 -62
rect 247 -73 251 -58
rect 273 -73 277 -50
rect 364 -54 368 -37
rect 390 -52 394 -37
rect 445 -52 449 -11
rect 693 -11 719 -9
rect 968 -9 1238 -7
rect 968 -11 1212 -9
rect 485 -23 493 -19
rect 497 -23 512 -19
rect 516 -23 530 -19
rect 534 -23 544 -19
rect 548 -23 745 -19
rect 749 -23 764 -19
rect 768 -23 782 -19
rect 786 -23 796 -19
rect 800 -23 862 -19
rect 866 -23 881 -19
rect 885 -23 899 -19
rect 903 -23 913 -19
rect 917 -21 933 -19
rect 937 -21 939 -19
rect 917 -23 939 -21
rect 488 -33 492 -23
rect 518 -33 522 -23
rect 530 -33 534 -23
rect 740 -33 744 -23
rect 770 -33 774 -23
rect 782 -33 786 -23
rect 857 -33 861 -23
rect 899 -33 903 -23
rect 503 -46 507 -37
rect 503 -50 522 -46
rect 348 -58 380 -54
rect 390 -56 449 -52
rect 518 -54 522 -50
rect 544 -52 548 -37
rect 755 -46 759 -37
rect 796 -46 800 -37
rect 707 -50 747 -46
rect 755 -50 774 -46
rect 330 -66 337 -62
rect 348 -73 352 -58
rect 390 -73 394 -56
rect 518 -58 534 -54
rect 544 -56 550 -52
rect 743 -54 747 -50
rect 770 -54 774 -50
rect 796 -50 876 -46
rect 518 -73 522 -58
rect 544 -73 548 -56
rect 743 -58 758 -54
rect 770 -58 786 -54
rect 695 -66 743 -62
rect 770 -73 774 -58
rect 796 -73 800 -50
rect 887 -54 891 -37
rect 913 -52 917 -37
rect 968 -52 972 -11
rect 1216 -11 1242 -9
rect 1008 -23 1016 -19
rect 1020 -23 1035 -19
rect 1039 -23 1053 -19
rect 1057 -23 1067 -19
rect 1071 -23 1268 -19
rect 1272 -23 1287 -19
rect 1291 -23 1305 -19
rect 1309 -23 1319 -19
rect 1323 -23 1385 -19
rect 1389 -23 1404 -19
rect 1408 -23 1422 -19
rect 1426 -23 1436 -19
rect 1440 -21 1456 -19
rect 1460 -21 1462 -19
rect 1440 -23 1462 -21
rect 1011 -33 1015 -23
rect 1041 -33 1045 -23
rect 1053 -33 1057 -23
rect 1263 -33 1267 -23
rect 1293 -33 1297 -23
rect 1305 -33 1309 -23
rect 1380 -33 1384 -23
rect 1422 -33 1426 -23
rect 1026 -46 1030 -37
rect 1026 -50 1045 -46
rect 871 -58 903 -54
rect 913 -56 972 -52
rect 1041 -54 1045 -50
rect 1067 -52 1071 -37
rect 1278 -46 1282 -37
rect 1319 -46 1323 -37
rect 1230 -50 1270 -46
rect 1278 -50 1297 -46
rect 853 -66 860 -62
rect 871 -73 875 -58
rect 913 -73 917 -56
rect 1041 -58 1057 -54
rect 1067 -56 1073 -52
rect 1266 -54 1270 -50
rect 1293 -54 1297 -50
rect 1319 -50 1399 -46
rect 1041 -73 1045 -58
rect 1067 -73 1071 -56
rect 1266 -58 1281 -54
rect 1293 -58 1309 -54
rect 1218 -66 1266 -62
rect 1293 -73 1297 -58
rect 1319 -73 1323 -50
rect 1410 -54 1414 -37
rect 1436 -52 1440 -37
rect 1394 -58 1426 -54
rect 1436 -56 1480 -52
rect 1376 -66 1383 -62
rect 1394 -73 1398 -58
rect 1436 -73 1440 -56
rect -558 -85 -554 -77
rect -516 -85 -512 -77
rect -306 -85 -302 -77
rect -264 -85 -260 -77
rect -189 -85 -185 -77
rect -159 -85 -155 -77
rect -147 -85 -143 -77
rect -612 -89 -553 -85
rect -549 -89 -532 -85
rect -528 -89 -516 -85
rect -512 -89 -501 -85
rect -497 -89 -301 -85
rect -297 -89 -280 -85
rect -276 -89 -264 -85
rect -260 -89 -249 -85
rect -245 -89 -184 -85
rect -180 -89 -163 -85
rect -159 -89 -147 -85
rect -143 -89 -132 -85
rect -128 -87 -121 -85
rect -35 -85 -31 -77
rect 7 -85 11 -77
rect 217 -85 221 -77
rect 259 -85 263 -77
rect 334 -85 338 -77
rect 364 -85 368 -77
rect 376 -85 380 -77
rect -117 -87 -30 -85
rect -128 -89 -30 -87
rect -26 -89 -9 -85
rect -5 -89 7 -85
rect 11 -89 22 -85
rect 26 -89 222 -85
rect 226 -89 243 -85
rect 247 -89 259 -85
rect 263 -89 274 -85
rect 278 -89 339 -85
rect 343 -89 360 -85
rect 364 -89 376 -85
rect 380 -89 391 -85
rect 395 -87 402 -85
rect 488 -85 492 -77
rect 530 -85 534 -77
rect 740 -85 744 -77
rect 782 -85 786 -77
rect 857 -85 861 -77
rect 887 -85 891 -77
rect 899 -85 903 -77
rect 406 -87 493 -85
rect 395 -89 493 -87
rect 497 -89 514 -85
rect 518 -89 530 -85
rect 534 -89 545 -85
rect 549 -89 745 -85
rect 749 -89 766 -85
rect 770 -89 782 -85
rect 786 -89 797 -85
rect 801 -89 862 -85
rect 866 -89 883 -85
rect 887 -89 899 -85
rect 903 -89 914 -85
rect 918 -87 925 -85
rect 1011 -85 1015 -77
rect 1053 -85 1057 -77
rect 1263 -85 1267 -77
rect 1305 -85 1309 -77
rect 1380 -85 1384 -77
rect 1410 -85 1414 -77
rect 1422 -85 1426 -77
rect 929 -87 1016 -85
rect 918 -89 1016 -87
rect 1020 -89 1037 -85
rect 1041 -89 1053 -85
rect 1057 -89 1068 -85
rect 1072 -89 1268 -85
rect 1272 -89 1289 -85
rect 1293 -89 1305 -85
rect 1309 -89 1320 -85
rect 1324 -89 1385 -85
rect 1389 -89 1406 -85
rect 1410 -89 1422 -85
rect 1426 -89 1437 -85
rect 1441 -87 1448 -85
rect 1452 -87 1480 -85
rect 1441 -89 1480 -87
<< metal2 >>
rect -504 115 -500 148
rect -269 115 -265 148
rect -502 111 -492 115
rect -267 111 -257 115
rect -496 71 -492 111
rect -496 67 -477 71
rect -500 45 -490 49
rect -494 7 -490 45
rect -434 7 -430 88
rect -261 71 -257 111
rect -261 67 -242 71
rect -410 49 -408 53
rect -410 7 -406 49
rect -265 45 -255 49
rect -259 7 -255 45
rect -199 7 -195 88
rect -175 49 -173 53
rect -175 7 -171 49
rect -121 -83 -117 -1
rect -113 -17 -109 148
rect 19 115 23 148
rect 254 115 258 148
rect 21 111 31 115
rect 256 111 266 115
rect 27 71 31 111
rect 27 67 46 71
rect 23 45 33 49
rect 29 7 33 45
rect 89 7 93 88
rect 262 71 266 111
rect 262 67 281 71
rect 113 49 115 53
rect 113 7 117 49
rect 258 45 268 49
rect 264 7 268 45
rect 324 7 328 88
rect 348 49 350 53
rect 348 7 352 49
rect 402 -83 406 -1
rect 410 -17 414 148
rect 542 115 546 148
rect 777 115 781 148
rect 544 111 554 115
rect 779 111 789 115
rect 550 71 554 111
rect 550 67 569 71
rect 546 45 556 49
rect 552 7 556 45
rect 612 7 616 88
rect 785 71 789 111
rect 785 67 804 71
rect 636 49 638 53
rect 636 7 640 49
rect 781 45 791 49
rect 787 7 791 45
rect 847 7 851 88
rect 871 49 873 53
rect 871 7 875 49
rect 925 -83 929 -1
rect 933 -17 937 148
rect 1065 115 1069 148
rect 1300 115 1304 148
rect 1067 111 1077 115
rect 1302 111 1312 115
rect 1073 71 1077 111
rect 1073 67 1092 71
rect 1069 45 1079 49
rect 1075 7 1079 45
rect 1135 7 1139 88
rect 1308 71 1312 111
rect 1308 67 1327 71
rect 1159 49 1161 53
rect 1159 7 1163 49
rect 1304 45 1314 49
rect 1310 7 1314 45
rect 1370 7 1374 88
rect 1394 49 1396 53
rect 1394 7 1398 49
rect 1448 -83 1452 -1
rect 1456 -17 1460 148
<< ntransistor >>
rect -464 94 -461 102
rect -449 94 -446 102
rect -531 55 -528 63
rect -516 55 -513 63
rect -396 59 -393 67
rect -381 59 -378 67
rect -464 11 -461 19
rect -449 11 -446 19
rect -550 -79 -547 -71
rect -535 -79 -532 -71
rect -508 -79 -506 -71
rect -229 94 -226 102
rect -214 94 -211 102
rect -296 55 -293 63
rect -281 55 -278 63
rect -161 59 -158 67
rect -146 59 -143 67
rect -229 11 -226 19
rect -214 11 -211 19
rect -298 -79 -295 -71
rect -283 -79 -280 -71
rect -256 -79 -254 -71
rect -181 -79 -178 -71
rect -166 -79 -163 -71
rect -139 -79 -137 -71
rect 59 94 62 102
rect 74 94 77 102
rect -8 55 -5 63
rect 7 55 10 63
rect 127 59 130 67
rect 142 59 145 67
rect 59 11 62 19
rect 74 11 77 19
rect -27 -79 -24 -71
rect -12 -79 -9 -71
rect 15 -79 17 -71
rect 294 94 297 102
rect 309 94 312 102
rect 227 55 230 63
rect 242 55 245 63
rect 362 59 365 67
rect 377 59 380 67
rect 294 11 297 19
rect 309 11 312 19
rect 225 -79 228 -71
rect 240 -79 243 -71
rect 267 -79 269 -71
rect 342 -79 345 -71
rect 357 -79 360 -71
rect 384 -79 386 -71
rect 582 94 585 102
rect 597 94 600 102
rect 515 55 518 63
rect 530 55 533 63
rect 650 59 653 67
rect 665 59 668 67
rect 582 11 585 19
rect 597 11 600 19
rect 496 -79 499 -71
rect 511 -79 514 -71
rect 538 -79 540 -71
rect 817 94 820 102
rect 832 94 835 102
rect 750 55 753 63
rect 765 55 768 63
rect 885 59 888 67
rect 900 59 903 67
rect 817 11 820 19
rect 832 11 835 19
rect 748 -79 751 -71
rect 763 -79 766 -71
rect 790 -79 792 -71
rect 865 -79 868 -71
rect 880 -79 883 -71
rect 907 -79 909 -71
rect 1105 94 1108 102
rect 1120 94 1123 102
rect 1038 55 1041 63
rect 1053 55 1056 63
rect 1173 59 1176 67
rect 1188 59 1191 67
rect 1105 11 1108 19
rect 1120 11 1123 19
rect 1019 -79 1022 -71
rect 1034 -79 1037 -71
rect 1061 -79 1063 -71
rect 1340 94 1343 102
rect 1355 94 1358 102
rect 1273 55 1276 63
rect 1288 55 1291 63
rect 1408 59 1411 67
rect 1423 59 1426 67
rect 1340 11 1343 19
rect 1355 11 1358 19
rect 1271 -79 1274 -71
rect 1286 -79 1289 -71
rect 1313 -79 1315 -71
rect 1388 -79 1391 -71
rect 1403 -79 1406 -71
rect 1430 -79 1432 -71
<< ptransistor >>
rect -464 134 -461 142
rect -449 134 -446 142
rect -229 134 -226 142
rect -214 134 -211 142
rect -531 95 -528 103
rect -516 95 -513 103
rect -396 99 -393 107
rect -381 99 -378 107
rect -296 95 -293 103
rect -281 95 -278 103
rect -464 51 -461 59
rect -449 51 -446 59
rect -550 -39 -547 -31
rect -535 -39 -532 -31
rect -508 -39 -506 -31
rect -161 99 -158 107
rect -146 99 -143 107
rect -229 51 -226 59
rect -214 51 -211 59
rect -298 -39 -295 -31
rect -283 -39 -280 -31
rect -256 -39 -254 -31
rect -181 -39 -178 -31
rect -166 -39 -163 -31
rect -139 -39 -137 -31
rect 59 134 62 142
rect 74 134 77 142
rect 294 134 297 142
rect 309 134 312 142
rect -8 95 -5 103
rect 7 95 10 103
rect 127 99 130 107
rect 142 99 145 107
rect 227 95 230 103
rect 242 95 245 103
rect 59 51 62 59
rect 74 51 77 59
rect -27 -39 -24 -31
rect -12 -39 -9 -31
rect 15 -39 17 -31
rect 362 99 365 107
rect 377 99 380 107
rect 294 51 297 59
rect 309 51 312 59
rect 225 -39 228 -31
rect 240 -39 243 -31
rect 267 -39 269 -31
rect 342 -39 345 -31
rect 357 -39 360 -31
rect 384 -39 386 -31
rect 582 134 585 142
rect 597 134 600 142
rect 817 134 820 142
rect 832 134 835 142
rect 515 95 518 103
rect 530 95 533 103
rect 650 99 653 107
rect 665 99 668 107
rect 750 95 753 103
rect 765 95 768 103
rect 582 51 585 59
rect 597 51 600 59
rect 496 -39 499 -31
rect 511 -39 514 -31
rect 538 -39 540 -31
rect 885 99 888 107
rect 900 99 903 107
rect 817 51 820 59
rect 832 51 835 59
rect 748 -39 751 -31
rect 763 -39 766 -31
rect 790 -39 792 -31
rect 865 -39 868 -31
rect 880 -39 883 -31
rect 907 -39 909 -31
rect 1105 134 1108 142
rect 1120 134 1123 142
rect 1340 134 1343 142
rect 1355 134 1358 142
rect 1038 95 1041 103
rect 1053 95 1056 103
rect 1173 99 1176 107
rect 1188 99 1191 107
rect 1273 95 1276 103
rect 1288 95 1291 103
rect 1105 51 1108 59
rect 1120 51 1123 59
rect 1019 -39 1022 -31
rect 1034 -39 1037 -31
rect 1061 -39 1063 -31
rect 1408 99 1411 107
rect 1423 99 1426 107
rect 1340 51 1343 59
rect 1355 51 1358 59
rect 1271 -39 1274 -31
rect 1286 -39 1289 -31
rect 1313 -39 1315 -31
rect 1388 -39 1391 -31
rect 1403 -39 1406 -31
rect 1430 -39 1432 -31
<< polycontact >>
rect -454 115 -450 119
rect -469 107 -465 111
rect -219 115 -215 119
rect -234 107 -230 111
rect -590 78 -586 82
rect -598 70 -594 74
rect -564 78 -560 82
rect -521 76 -517 80
rect -386 80 -382 84
rect -564 66 -560 70
rect -536 68 -532 72
rect -401 72 -397 76
rect -345 78 -341 82
rect -454 32 -450 36
rect -469 24 -465 28
rect -357 -13 -353 -9
rect -512 -58 -508 -54
rect -496 -56 -492 -52
rect -286 76 -282 80
rect -151 80 -147 84
rect -331 66 -327 70
rect -301 68 -297 72
rect -166 72 -162 76
rect -104 78 -100 82
rect -219 32 -215 36
rect -234 24 -230 28
rect -331 -9 -327 -5
rect -343 -50 -339 -46
rect -288 -58 -284 -54
rect -260 -58 -256 -54
rect -355 -66 -351 -62
rect -303 -66 -299 -62
rect -170 -50 -166 -46
rect -186 -66 -182 -62
rect -143 -58 -139 -54
rect 69 115 73 119
rect 54 107 58 111
rect 304 115 308 119
rect 289 107 293 111
rect -67 78 -63 82
rect -75 70 -71 74
rect -41 78 -37 82
rect 2 76 6 80
rect 137 80 141 84
rect -41 66 -37 70
rect -13 68 -9 72
rect 122 72 126 76
rect 178 78 182 82
rect 69 32 73 36
rect 54 24 58 28
rect 166 -13 170 -9
rect 11 -58 15 -54
rect 27 -56 31 -52
rect 237 76 241 80
rect 372 80 376 84
rect 192 66 196 70
rect 222 68 226 72
rect 357 72 361 76
rect 419 78 423 82
rect 304 32 308 36
rect 289 24 293 28
rect 192 -9 196 -5
rect 180 -50 184 -46
rect 235 -58 239 -54
rect 263 -58 267 -54
rect 168 -66 172 -62
rect 220 -66 224 -62
rect 353 -50 357 -46
rect 337 -66 341 -62
rect 380 -58 384 -54
rect 592 115 596 119
rect 577 107 581 111
rect 827 115 831 119
rect 812 107 816 111
rect 456 78 460 82
rect 448 70 452 74
rect 482 78 486 82
rect 525 76 529 80
rect 660 80 664 84
rect 482 66 486 70
rect 510 68 514 72
rect 645 72 649 76
rect 701 78 705 82
rect 592 32 596 36
rect 577 24 581 28
rect 689 -13 693 -9
rect 534 -58 538 -54
rect 550 -56 554 -52
rect 760 76 764 80
rect 895 80 899 84
rect 715 66 719 70
rect 745 68 749 72
rect 880 72 884 76
rect 942 78 946 82
rect 827 32 831 36
rect 812 24 816 28
rect 715 -9 719 -5
rect 703 -50 707 -46
rect 758 -58 762 -54
rect 786 -58 790 -54
rect 691 -66 695 -62
rect 743 -66 747 -62
rect 876 -50 880 -46
rect 860 -66 864 -62
rect 903 -58 907 -54
rect 1115 115 1119 119
rect 1100 107 1104 111
rect 1350 115 1354 119
rect 1335 107 1339 111
rect 979 78 983 82
rect 971 70 975 74
rect 1005 78 1009 82
rect 1048 76 1052 80
rect 1183 80 1187 84
rect 1005 66 1009 70
rect 1033 68 1037 72
rect 1168 72 1172 76
rect 1224 78 1228 82
rect 1115 32 1119 36
rect 1100 24 1104 28
rect 1212 -13 1216 -9
rect 1057 -58 1061 -54
rect 1073 -56 1077 -52
rect 1283 76 1287 80
rect 1418 80 1422 84
rect 1238 66 1242 70
rect 1268 68 1272 72
rect 1403 72 1407 76
rect 1465 78 1469 82
rect 1350 32 1354 36
rect 1335 24 1339 28
rect 1238 -9 1242 -5
rect 1226 -50 1230 -46
rect 1281 -58 1285 -54
rect 1309 -58 1313 -54
rect 1214 -66 1218 -62
rect 1266 -66 1270 -62
rect 1399 -50 1403 -46
rect 1383 -66 1387 -62
rect 1426 -58 1430 -54
<< ndcontact >>
rect -472 96 -468 100
rect -442 96 -438 100
rect -237 96 -233 100
rect -539 57 -535 61
rect -509 57 -505 61
rect -404 61 -400 65
rect -374 61 -370 65
rect -472 13 -468 17
rect -442 13 -438 17
rect -558 -77 -554 -73
rect -528 -77 -524 -73
rect -516 -77 -512 -73
rect -502 -77 -498 -73
rect -207 96 -203 100
rect -304 57 -300 61
rect -274 57 -270 61
rect -169 61 -165 65
rect -139 61 -135 65
rect -237 13 -233 17
rect -207 13 -203 17
rect -306 -77 -302 -73
rect -276 -77 -272 -73
rect -264 -77 -260 -73
rect -250 -77 -246 -73
rect -189 -77 -185 -73
rect -175 -77 -171 -73
rect -159 -77 -155 -73
rect -147 -77 -143 -73
rect -133 -77 -129 -73
rect 51 96 55 100
rect 81 96 85 100
rect 286 96 290 100
rect -16 57 -12 61
rect 14 57 18 61
rect 119 61 123 65
rect 149 61 153 65
rect 51 13 55 17
rect 81 13 85 17
rect -35 -77 -31 -73
rect -5 -77 -1 -73
rect 7 -77 11 -73
rect 21 -77 25 -73
rect 316 96 320 100
rect 219 57 223 61
rect 249 57 253 61
rect 354 61 358 65
rect 384 61 388 65
rect 286 13 290 17
rect 316 13 320 17
rect 217 -77 221 -73
rect 247 -77 251 -73
rect 259 -77 263 -73
rect 273 -77 277 -73
rect 334 -77 338 -73
rect 348 -77 352 -73
rect 364 -77 368 -73
rect 376 -77 380 -73
rect 390 -77 394 -73
rect 574 96 578 100
rect 604 96 608 100
rect 809 96 813 100
rect 507 57 511 61
rect 537 57 541 61
rect 642 61 646 65
rect 672 61 676 65
rect 574 13 578 17
rect 604 13 608 17
rect 488 -77 492 -73
rect 518 -77 522 -73
rect 530 -77 534 -73
rect 544 -77 548 -73
rect 839 96 843 100
rect 742 57 746 61
rect 772 57 776 61
rect 877 61 881 65
rect 907 61 911 65
rect 809 13 813 17
rect 839 13 843 17
rect 740 -77 744 -73
rect 770 -77 774 -73
rect 782 -77 786 -73
rect 796 -77 800 -73
rect 857 -77 861 -73
rect 871 -77 875 -73
rect 887 -77 891 -73
rect 899 -77 903 -73
rect 913 -77 917 -73
rect 1097 96 1101 100
rect 1127 96 1131 100
rect 1332 96 1336 100
rect 1030 57 1034 61
rect 1060 57 1064 61
rect 1165 61 1169 65
rect 1195 61 1199 65
rect 1097 13 1101 17
rect 1127 13 1131 17
rect 1011 -77 1015 -73
rect 1041 -77 1045 -73
rect 1053 -77 1057 -73
rect 1067 -77 1071 -73
rect 1362 96 1366 100
rect 1265 57 1269 61
rect 1295 57 1299 61
rect 1400 61 1404 65
rect 1430 61 1434 65
rect 1332 13 1336 17
rect 1362 13 1366 17
rect 1263 -77 1267 -73
rect 1293 -77 1297 -73
rect 1305 -77 1309 -73
rect 1319 -77 1323 -73
rect 1380 -77 1384 -73
rect 1394 -77 1398 -73
rect 1410 -77 1414 -73
rect 1422 -77 1426 -73
rect 1436 -77 1440 -73
<< pdcontact >>
rect -472 136 -468 140
rect -457 136 -453 140
rect -442 136 -438 140
rect -237 136 -233 140
rect -222 136 -218 140
rect -207 136 -203 140
rect -539 97 -535 101
rect -524 97 -520 101
rect -509 97 -505 101
rect -404 101 -400 105
rect -389 101 -385 105
rect -374 101 -370 105
rect -304 97 -300 101
rect -289 97 -285 101
rect -274 97 -270 101
rect -472 53 -468 57
rect -457 53 -453 57
rect -442 53 -438 57
rect -558 -37 -554 -33
rect -543 -37 -539 -33
rect -528 -37 -524 -33
rect -516 -37 -512 -33
rect -502 -37 -498 -33
rect -169 101 -165 105
rect -154 101 -150 105
rect -139 101 -135 105
rect -237 53 -233 57
rect -222 53 -218 57
rect -207 53 -203 57
rect -306 -37 -302 -33
rect -291 -37 -287 -33
rect -276 -37 -272 -33
rect -264 -37 -260 -33
rect -250 -37 -246 -33
rect -189 -37 -185 -33
rect -159 -37 -155 -33
rect -147 -37 -143 -33
rect -133 -37 -129 -33
rect 51 136 55 140
rect 66 136 70 140
rect 81 136 85 140
rect 286 136 290 140
rect 301 136 305 140
rect 316 136 320 140
rect -16 97 -12 101
rect -1 97 3 101
rect 14 97 18 101
rect 119 101 123 105
rect 134 101 138 105
rect 149 101 153 105
rect 219 97 223 101
rect 234 97 238 101
rect 249 97 253 101
rect 51 53 55 57
rect 66 53 70 57
rect 81 53 85 57
rect -35 -37 -31 -33
rect -20 -37 -16 -33
rect -5 -37 -1 -33
rect 7 -37 11 -33
rect 21 -37 25 -33
rect 354 101 358 105
rect 369 101 373 105
rect 384 101 388 105
rect 286 53 290 57
rect 301 53 305 57
rect 316 53 320 57
rect 217 -37 221 -33
rect 232 -37 236 -33
rect 247 -37 251 -33
rect 259 -37 263 -33
rect 273 -37 277 -33
rect 334 -37 338 -33
rect 364 -37 368 -33
rect 376 -37 380 -33
rect 390 -37 394 -33
rect 574 136 578 140
rect 589 136 593 140
rect 604 136 608 140
rect 809 136 813 140
rect 824 136 828 140
rect 839 136 843 140
rect 507 97 511 101
rect 522 97 526 101
rect 537 97 541 101
rect 642 101 646 105
rect 657 101 661 105
rect 672 101 676 105
rect 742 97 746 101
rect 757 97 761 101
rect 772 97 776 101
rect 574 53 578 57
rect 589 53 593 57
rect 604 53 608 57
rect 488 -37 492 -33
rect 503 -37 507 -33
rect 518 -37 522 -33
rect 530 -37 534 -33
rect 544 -37 548 -33
rect 877 101 881 105
rect 892 101 896 105
rect 907 101 911 105
rect 809 53 813 57
rect 824 53 828 57
rect 839 53 843 57
rect 740 -37 744 -33
rect 755 -37 759 -33
rect 770 -37 774 -33
rect 782 -37 786 -33
rect 796 -37 800 -33
rect 857 -37 861 -33
rect 887 -37 891 -33
rect 899 -37 903 -33
rect 913 -37 917 -33
rect 1097 136 1101 140
rect 1112 136 1116 140
rect 1127 136 1131 140
rect 1332 136 1336 140
rect 1347 136 1351 140
rect 1362 136 1366 140
rect 1030 97 1034 101
rect 1045 97 1049 101
rect 1060 97 1064 101
rect 1165 101 1169 105
rect 1180 101 1184 105
rect 1195 101 1199 105
rect 1265 97 1269 101
rect 1280 97 1284 101
rect 1295 97 1299 101
rect 1097 53 1101 57
rect 1112 53 1116 57
rect 1127 53 1131 57
rect 1011 -37 1015 -33
rect 1026 -37 1030 -33
rect 1041 -37 1045 -33
rect 1053 -37 1057 -33
rect 1067 -37 1071 -33
rect 1400 101 1404 105
rect 1415 101 1419 105
rect 1430 101 1434 105
rect 1332 53 1336 57
rect 1347 53 1351 57
rect 1362 53 1366 57
rect 1263 -37 1267 -33
rect 1278 -37 1282 -33
rect 1293 -37 1297 -33
rect 1305 -37 1309 -33
rect 1319 -37 1323 -33
rect 1380 -37 1384 -33
rect 1410 -37 1414 -33
rect 1422 -37 1426 -33
rect 1436 -37 1440 -33
<< nbccdiffcontact >>
rect -516 -23 -512 -19
rect -264 -23 -260 -19
rect -147 -23 -143 -19
rect 7 -23 11 -19
rect 259 -23 263 -19
rect 376 -23 380 -19
rect 530 -23 534 -19
rect 782 -23 786 -19
rect 899 -23 903 -19
rect 1053 -23 1057 -19
rect 1305 -23 1309 -19
rect 1422 -23 1426 -19
<< m2contact >>
rect -504 148 -500 152
rect -269 148 -265 152
rect -113 148 -109 152
rect 19 148 23 152
rect 254 148 258 152
rect 410 148 414 152
rect 542 148 546 152
rect 777 148 781 152
rect 933 148 937 152
rect 1065 148 1069 152
rect 1300 148 1304 152
rect 1456 148 1460 152
rect -506 111 -502 115
rect -438 84 -434 88
rect -271 111 -267 115
rect -504 45 -500 49
rect -477 67 -473 71
rect -203 84 -199 88
rect -408 49 -404 53
rect -269 45 -265 49
rect -242 67 -238 71
rect 17 111 21 115
rect 85 84 89 88
rect 252 111 256 115
rect -173 49 -169 53
rect 19 45 23 49
rect 46 67 50 71
rect 320 84 324 88
rect 115 49 119 53
rect 254 45 258 49
rect 281 67 285 71
rect 540 111 544 115
rect 608 84 612 88
rect 775 111 779 115
rect 350 49 354 53
rect 542 45 546 49
rect 569 67 573 71
rect 843 84 847 88
rect 638 49 642 53
rect 777 45 781 49
rect 804 67 808 71
rect 1063 111 1067 115
rect 1131 84 1135 88
rect 1298 111 1302 115
rect 873 49 877 53
rect 1065 45 1069 49
rect 1092 67 1096 71
rect 1366 84 1370 88
rect 1161 49 1165 53
rect 1300 45 1304 49
rect 1327 67 1331 71
rect 1396 49 1400 53
rect -494 3 -490 7
rect -434 3 -430 7
rect -410 3 -406 7
rect -259 3 -255 7
rect -199 3 -195 7
rect -175 3 -171 7
rect -121 -1 -117 3
rect 29 3 33 7
rect 89 3 93 7
rect 113 3 117 7
rect 264 3 268 7
rect 324 3 328 7
rect 348 3 352 7
rect 402 -1 406 3
rect 552 3 556 7
rect 612 3 616 7
rect 636 3 640 7
rect 787 3 791 7
rect 847 3 851 7
rect 871 3 875 7
rect 925 -1 929 3
rect 1075 3 1079 7
rect 1135 3 1139 7
rect 1159 3 1163 7
rect 1310 3 1314 7
rect 1370 3 1374 7
rect 1394 3 1398 7
rect 1448 -1 1452 3
rect -113 -21 -109 -17
rect 410 -21 414 -17
rect 933 -21 937 -17
rect 1456 -21 1460 -17
rect -121 -87 -117 -83
rect 402 -87 406 -83
rect 925 -87 929 -83
rect 1448 -87 1452 -83
<< psubstratepcontact >>
rect -467 84 -463 88
rect -446 84 -442 88
rect -534 45 -530 49
rect -513 45 -509 49
rect -399 49 -395 53
rect -378 49 -374 53
rect -467 1 -463 5
rect -446 1 -442 5
rect -553 -89 -549 -85
rect -532 -89 -528 -85
rect -516 -89 -512 -85
rect -501 -89 -497 -85
rect -232 84 -228 88
rect -211 84 -207 88
rect -299 45 -295 49
rect -278 45 -274 49
rect -164 49 -160 53
rect -143 49 -139 53
rect -232 1 -228 5
rect -211 1 -207 5
rect -301 -89 -297 -85
rect -280 -89 -276 -85
rect -264 -89 -260 -85
rect -249 -89 -245 -85
rect -184 -89 -180 -85
rect -163 -89 -159 -85
rect -147 -89 -143 -85
rect -132 -89 -128 -85
rect 56 84 60 88
rect 77 84 81 88
rect -11 45 -7 49
rect 10 45 14 49
rect 124 49 128 53
rect 145 49 149 53
rect 56 1 60 5
rect 77 1 81 5
rect -30 -89 -26 -85
rect -9 -89 -5 -85
rect 7 -89 11 -85
rect 22 -89 26 -85
rect 291 84 295 88
rect 312 84 316 88
rect 224 45 228 49
rect 245 45 249 49
rect 359 49 363 53
rect 380 49 384 53
rect 291 1 295 5
rect 312 1 316 5
rect 222 -89 226 -85
rect 243 -89 247 -85
rect 259 -89 263 -85
rect 274 -89 278 -85
rect 339 -89 343 -85
rect 360 -89 364 -85
rect 376 -89 380 -85
rect 391 -89 395 -85
rect 579 84 583 88
rect 600 84 604 88
rect 512 45 516 49
rect 533 45 537 49
rect 647 49 651 53
rect 668 49 672 53
rect 579 1 583 5
rect 600 1 604 5
rect 493 -89 497 -85
rect 514 -89 518 -85
rect 530 -89 534 -85
rect 545 -89 549 -85
rect 814 84 818 88
rect 835 84 839 88
rect 747 45 751 49
rect 768 45 772 49
rect 882 49 886 53
rect 903 49 907 53
rect 814 1 818 5
rect 835 1 839 5
rect 745 -89 749 -85
rect 766 -89 770 -85
rect 782 -89 786 -85
rect 797 -89 801 -85
rect 862 -89 866 -85
rect 883 -89 887 -85
rect 899 -89 903 -85
rect 914 -89 918 -85
rect 1102 84 1106 88
rect 1123 84 1127 88
rect 1035 45 1039 49
rect 1056 45 1060 49
rect 1170 49 1174 53
rect 1191 49 1195 53
rect 1102 1 1106 5
rect 1123 1 1127 5
rect 1016 -89 1020 -85
rect 1037 -89 1041 -85
rect 1053 -89 1057 -85
rect 1068 -89 1072 -85
rect 1337 84 1341 88
rect 1358 84 1362 88
rect 1270 45 1274 49
rect 1291 45 1295 49
rect 1405 49 1409 53
rect 1426 49 1430 53
rect 1337 1 1341 5
rect 1358 1 1362 5
rect 1268 -89 1272 -85
rect 1289 -89 1293 -85
rect 1305 -89 1309 -85
rect 1320 -89 1324 -85
rect 1385 -89 1389 -85
rect 1406 -89 1410 -85
rect 1422 -89 1426 -85
rect 1437 -89 1441 -85
<< nsubstratencontact >>
rect -467 150 -463 154
rect -448 150 -444 154
rect -232 150 -228 154
rect -213 150 -209 154
rect -534 111 -530 115
rect -515 111 -511 115
rect -399 115 -395 119
rect -380 115 -376 119
rect -299 111 -295 115
rect -280 111 -276 115
rect -164 115 -160 119
rect -145 115 -141 119
rect -467 67 -463 71
rect -448 67 -444 71
rect -553 -23 -549 -19
rect -534 -23 -530 -19
rect -502 -23 -498 -19
rect -232 67 -228 71
rect -213 67 -209 71
rect -301 -23 -297 -19
rect -282 -23 -278 -19
rect -250 -23 -246 -19
rect -184 -23 -180 -19
rect -165 -23 -161 -19
rect -133 -23 -129 -19
rect 56 150 60 154
rect 75 150 79 154
rect 291 150 295 154
rect 310 150 314 154
rect -11 111 -7 115
rect 8 111 12 115
rect 124 115 128 119
rect 143 115 147 119
rect 224 111 228 115
rect 243 111 247 115
rect 359 115 363 119
rect 378 115 382 119
rect 56 67 60 71
rect 75 67 79 71
rect -30 -23 -26 -19
rect -11 -23 -7 -19
rect 21 -23 25 -19
rect 291 67 295 71
rect 310 67 314 71
rect 222 -23 226 -19
rect 241 -23 245 -19
rect 273 -23 277 -19
rect 339 -23 343 -19
rect 358 -23 362 -19
rect 390 -23 394 -19
rect 579 150 583 154
rect 598 150 602 154
rect 814 150 818 154
rect 833 150 837 154
rect 512 111 516 115
rect 531 111 535 115
rect 647 115 651 119
rect 666 115 670 119
rect 747 111 751 115
rect 766 111 770 115
rect 882 115 886 119
rect 901 115 905 119
rect 579 67 583 71
rect 598 67 602 71
rect 493 -23 497 -19
rect 512 -23 516 -19
rect 544 -23 548 -19
rect 814 67 818 71
rect 833 67 837 71
rect 745 -23 749 -19
rect 764 -23 768 -19
rect 796 -23 800 -19
rect 862 -23 866 -19
rect 881 -23 885 -19
rect 913 -23 917 -19
rect 1102 150 1106 154
rect 1121 150 1125 154
rect 1337 150 1341 154
rect 1356 150 1360 154
rect 1035 111 1039 115
rect 1054 111 1058 115
rect 1170 115 1174 119
rect 1189 115 1193 119
rect 1270 111 1274 115
rect 1289 111 1293 115
rect 1405 115 1409 119
rect 1424 115 1428 119
rect 1102 67 1106 71
rect 1121 67 1125 71
rect 1016 -23 1020 -19
rect 1035 -23 1039 -19
rect 1067 -23 1071 -19
rect 1337 67 1341 71
rect 1356 67 1360 71
rect 1268 -23 1272 -19
rect 1287 -23 1291 -19
rect 1319 -23 1323 -19
rect 1385 -23 1389 -19
rect 1404 -23 1408 -19
rect 1436 -23 1440 -19
<< labels >>
rlabel metal1 -610 -54 -610 -54 3 ctrl
rlabel metal1 -39 151 -39 151 1 Vdd
rlabel metal1 -47 -87 -47 -87 1 gnd
rlabel polysilicon -596 163 -596 163 5 a0
rlabel polysilicon -588 163 -588 163 5 b0
rlabel polysilicon -73 162 -73 162 5 a1
rlabel polysilicon -65 162 -65 162 5 b1
rlabel polysilicon 450 161 450 161 5 a2
rlabel polysilicon 458 161 458 161 5 b2
rlabel polysilicon 973 161 973 161 5 a3
rlabel polysilicon 981 161 981 161 5 b3
rlabel metal1 1478 -54 1478 -54 7 Carry
rlabel polysilicon 1467 -102 1467 -102 1 s3
rlabel polysilicon 944 -101 944 -101 1 s2
rlabel polysilicon 421 -101 421 -101 1 s1
rlabel polysilicon -102 -101 -102 -101 1 s0
<< end >>
