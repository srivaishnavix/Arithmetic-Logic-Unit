* SPICE3 file created from DECODER.ext - technology: scmos


.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'

.option scale=1u

M1000 a_n57_n89# s0 gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1001 vdd a_n57_n5# a_156_n117# w_141_n119# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1002 vdd s1 a_150_111# w_135_109# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1003 d2 a_152_35# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1004 a_154_n41# s0 vdd w_139_n43# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1005 a_n57_n5# s1 gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1006 d1 a_154_n41# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1007 a_n57_n89# s0 vdd w_n70_n51# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1008 a_156_n157# a_n57_n89# gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1009 a_150_111# s1 a_150_71# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1010 a_152_35# a_n57_n89# vdd w_137_33# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1011 a_152_35# s1 a_152_n5# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1012 d1 a_154_n41# vdd w_139_n43# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1013 a_150_111# s0 vdd w_135_109# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1014 a_154_n41# a_n57_n5# a_154_n81# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1015 d3 a_150_111# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1016 a_156_n117# a_n57_n89# vdd w_141_n119# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1017 d2 a_152_35# vdd w_137_33# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1018 d0 a_156_n117# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1019 a_n57_n5# s1 vdd w_n70_33# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1020 vdd a_n57_n5# a_154_n41# w_139_n43# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1021 a_156_n117# a_n57_n5# a_156_n157# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1022 d3 a_150_111# vdd w_135_109# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1023 a_154_n81# s0 gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1024 a_150_71# s0 gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1025 d0 a_156_n117# vdd w_141_n119# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1026 a_152_n5# a_n57_n89# gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1027 vdd s1 a_152_35# w_137_33# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
C0 d0 0 11.468f 
C1 a_156_n117# 0 21.108f 
C2 d1 0 11.844f 
C3 a_154_n41# 0 21.108f 
C4 d2 0 12.22f 
C5 a_152_35# 0 21.108f 
C6 a_n57_n89# 0 0.121192p 
C7 gnd 0 0.1589p 
C8 a_n57_n5# 0 0.16038p 
C9 d3 0 12.596f 
C10 a_150_111# 0 21.108f 
C11 s1 0 0.179276p 
C12 s0 0 0.194784p 
C13 vdd 0 0.166212p 



Vs1 s1 gnd 0

Vs0 s0 gnd 0



.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(d3) v(d2)+2 v(d1)+4 v(d0)+6

.end
.endc