* SPICE3 file created from 4AND.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'

.option scale=1u

M1000 a_35_16# a1 Vdd w_20_14 CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1001 Vdd b1 a_35_16# w_20_14 CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1002 a_112_16# b2 a_112_n24# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1003 Vdd b0 a_n42_16# w_n57_14 CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1004 a_35_n24# a1 gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1005 a_n42_16# b0 a_n42_n24# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1006 Vdd b2 a_112_16# w_97_14 CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1007 a_189_16# a3 Vdd w_174_14 CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1008 s1 a_35_16# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1009 a_112_n24# a2 gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1010 s3 a_189_16# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1011 a_n42_16# a0 Vdd w_n57_14 CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1012 s0 a_n42_16# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1013 s1 a_35_16# Vdd w_20_14 CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1014 a_112_16# a2 Vdd w_97_14 CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1015 Vdd b3 a_189_16# w_174_14 CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1016 a_n42_n24# a0 gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1017 a_35_16# b1 a_35_n24# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1018 a_189_16# b3 a_189_n24# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1019 s2 a_112_16# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1020 s3 a_189_16# Vdd w_174_14 CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1021 s2 a_112_16# Vdd w_97_14 CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1022 a_189_n24# a3 gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1023 s0 a_n42_16# Vdd w_n57_14 CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
C0 gnd 0 50.572f 
C1 s3 0 23.720001f 
C2 s2 0 23.720001f 
C3 s1 0 23.720001f 
C4 s0 0 23.720001f 
C5 a_189_16# 0 21.108f 
C6 b3 0 20.639f 
C7 a_112_16# 0 21.108f 
C8 a3 0 20.639f 
C9 b2 0 20.639f 
C10 a_35_16# 0 21.108f 
C11 a2 0 20.639f 
C12 b1 0 20.639f 
C13 a_n42_16# 0 21.108f 
C14 a1 0 20.639f 
C15 b0 0 20.639f 
C16 a0 0 20.639f 
C17 Vdd 0 53.204f 

Va0 a0 gnd 0
Va1 a1 gnd 1
Va2 a2 gnd 0
Va3 a3 gnd 1

Vb0 b0 gnd 1
Vb1 b1 gnd 1
Vb2 b2 gnd 1
Vb3 b3 gnd 1



.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(a3) v(b3)+2 v(s3)+4 
plot v(a2) v(b2)+2 v(s2)+4 
plot v(a1) v(b1)+2 v(s1)+4 
plot v(a0) v(b0)+2 v(s0)+4 

.end
.endc