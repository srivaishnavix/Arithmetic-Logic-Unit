magic
tech scmos
timestamp 1701023198
<< nwell >>
rect -57 14 11 26
rect 20 14 88 26
rect 97 14 165 26
rect 174 14 242 26
<< polysilicon >>
rect -42 29 -39 58
rect -45 26 -39 29
rect -33 29 -30 58
rect 35 29 38 58
rect -33 26 -27 29
rect -45 24 -42 26
rect -30 24 -27 26
rect -3 24 -1 28
rect 32 26 38 29
rect 44 29 47 58
rect 112 29 115 58
rect 44 26 50 29
rect 32 24 35 26
rect 47 24 50 26
rect 74 24 76 28
rect 109 26 115 29
rect 121 29 124 58
rect 189 29 192 58
rect 121 26 127 29
rect 109 24 112 26
rect 124 24 127 26
rect 151 24 153 28
rect 186 26 192 29
rect 198 29 201 58
rect 198 26 204 29
rect 186 24 189 26
rect 201 24 204 26
rect 228 24 230 28
rect -45 -16 -42 16
rect -30 -16 -27 16
rect -3 -16 -1 16
rect 13 -1 15 3
rect -45 -26 -42 -24
rect -30 -26 -27 -24
rect -3 -26 -1 -24
rect 11 -49 15 -1
rect 32 -16 35 16
rect 47 -16 50 16
rect 74 -16 76 16
rect 90 -1 92 3
rect 32 -26 35 -24
rect 47 -26 50 -24
rect 74 -26 76 -24
rect 88 -49 92 -1
rect 109 -16 112 16
rect 124 -16 127 16
rect 151 -16 153 16
rect 167 -1 169 3
rect 109 -26 112 -24
rect 124 -26 127 -24
rect 151 -26 153 -24
rect 165 -49 169 -1
rect 186 -16 189 16
rect 201 -16 204 16
rect 228 -16 230 16
rect 244 -1 246 3
rect 186 -26 189 -24
rect 201 -26 204 -24
rect 228 -26 230 -24
rect 242 -49 246 -1
<< ndiffusion >>
rect -55 -18 -45 -16
rect -55 -22 -53 -18
rect -49 -22 -45 -18
rect -55 -24 -45 -22
rect -42 -24 -30 -16
rect -27 -18 -17 -16
rect -27 -22 -23 -18
rect -19 -22 -17 -18
rect -27 -24 -17 -22
rect -13 -18 -3 -16
rect -13 -22 -11 -18
rect -7 -22 -3 -18
rect -13 -24 -3 -22
rect -1 -18 9 -16
rect -1 -22 3 -18
rect 7 -22 9 -18
rect -1 -24 9 -22
rect 22 -18 32 -16
rect 22 -22 24 -18
rect 28 -22 32 -18
rect 22 -24 32 -22
rect 35 -24 47 -16
rect 50 -18 60 -16
rect 50 -22 54 -18
rect 58 -22 60 -18
rect 50 -24 60 -22
rect 64 -18 74 -16
rect 64 -22 66 -18
rect 70 -22 74 -18
rect 64 -24 74 -22
rect 76 -18 86 -16
rect 76 -22 80 -18
rect 84 -22 86 -18
rect 76 -24 86 -22
rect 99 -18 109 -16
rect 99 -22 101 -18
rect 105 -22 109 -18
rect 99 -24 109 -22
rect 112 -24 124 -16
rect 127 -18 137 -16
rect 127 -22 131 -18
rect 135 -22 137 -18
rect 127 -24 137 -22
rect 141 -18 151 -16
rect 141 -22 143 -18
rect 147 -22 151 -18
rect 141 -24 151 -22
rect 153 -18 163 -16
rect 153 -22 157 -18
rect 161 -22 163 -18
rect 153 -24 163 -22
rect 176 -18 186 -16
rect 176 -22 178 -18
rect 182 -22 186 -18
rect 176 -24 186 -22
rect 189 -24 201 -16
rect 204 -18 214 -16
rect 204 -22 208 -18
rect 212 -22 214 -18
rect 204 -24 214 -22
rect 218 -18 228 -16
rect 218 -22 220 -18
rect 224 -22 228 -18
rect 218 -24 228 -22
rect 230 -18 240 -16
rect 230 -22 234 -18
rect 238 -22 240 -18
rect 230 -24 240 -22
<< pdiffusion >>
rect -55 22 -45 24
rect -55 18 -53 22
rect -49 18 -45 22
rect -55 16 -45 18
rect -42 22 -30 24
rect -42 18 -38 22
rect -34 18 -30 22
rect -42 16 -30 18
rect -27 22 -17 24
rect -27 18 -23 22
rect -19 18 -17 22
rect -27 16 -17 18
rect -13 22 -3 24
rect -13 18 -11 22
rect -7 18 -3 22
rect -13 16 -3 18
rect -1 22 9 24
rect -1 18 3 22
rect 7 18 9 22
rect -1 16 9 18
rect 22 22 32 24
rect 22 18 24 22
rect 28 18 32 22
rect 22 16 32 18
rect 35 22 47 24
rect 35 18 39 22
rect 43 18 47 22
rect 35 16 47 18
rect 50 22 60 24
rect 50 18 54 22
rect 58 18 60 22
rect 50 16 60 18
rect 64 22 74 24
rect 64 18 66 22
rect 70 18 74 22
rect 64 16 74 18
rect 76 22 86 24
rect 76 18 80 22
rect 84 18 86 22
rect 76 16 86 18
rect 99 22 109 24
rect 99 18 101 22
rect 105 18 109 22
rect 99 16 109 18
rect 112 22 124 24
rect 112 18 116 22
rect 120 18 124 22
rect 112 16 124 18
rect 127 22 137 24
rect 127 18 131 22
rect 135 18 137 22
rect 127 16 137 18
rect 141 22 151 24
rect 141 18 143 22
rect 147 18 151 22
rect 141 16 151 18
rect 153 22 163 24
rect 153 18 157 22
rect 161 18 163 22
rect 153 16 163 18
rect 176 22 186 24
rect 176 18 178 22
rect 182 18 186 22
rect 176 16 186 18
rect 189 22 201 24
rect 189 18 193 22
rect 197 18 201 22
rect 189 16 201 18
rect 204 22 214 24
rect 204 18 208 22
rect 212 18 214 22
rect 204 16 214 18
rect 218 22 228 24
rect 218 18 220 22
rect 224 18 228 22
rect 218 16 228 18
rect 230 22 240 24
rect 230 18 234 22
rect 238 18 240 22
rect 230 16 240 18
<< metal1 >>
rect -57 32 -48 36
rect -44 32 -29 36
rect -25 32 -11 36
rect -7 32 3 36
rect 7 32 29 36
rect 33 32 48 36
rect 52 32 66 36
rect 70 32 80 36
rect 84 32 106 36
rect 110 32 125 36
rect 129 32 143 36
rect 147 32 157 36
rect 161 32 183 36
rect 187 32 202 36
rect 206 32 220 36
rect 224 32 234 36
rect 238 32 242 36
rect -53 22 -49 32
rect -23 22 -19 32
rect -11 22 -7 32
rect 24 22 28 32
rect 54 22 58 32
rect 66 22 70 32
rect 101 22 105 32
rect 131 22 135 32
rect 143 22 147 32
rect 178 22 182 32
rect 208 22 212 32
rect 220 22 224 32
rect -38 9 -34 18
rect -38 5 -19 9
rect -23 1 -19 5
rect 3 3 7 18
rect 39 9 43 18
rect 39 5 58 9
rect -23 -3 -7 1
rect 3 -1 9 3
rect 54 1 58 5
rect 80 3 84 18
rect 116 9 120 18
rect 116 5 135 9
rect -23 -18 -19 -3
rect 3 -18 7 -1
rect 54 -3 70 1
rect 80 -1 86 3
rect 131 1 135 5
rect 157 3 161 18
rect 193 9 197 18
rect 193 5 212 9
rect 54 -18 58 -3
rect 80 -18 84 -1
rect 131 -3 147 1
rect 157 -1 163 3
rect 208 1 212 5
rect 234 3 238 18
rect 131 -18 135 -3
rect 157 -18 161 -1
rect 208 -3 224 1
rect 234 -1 240 3
rect 208 -18 212 -3
rect 234 -18 238 -1
rect -53 -30 -49 -22
rect -11 -30 -7 -22
rect 24 -30 28 -22
rect 66 -30 70 -22
rect 101 -30 105 -22
rect 143 -30 147 -22
rect 178 -30 182 -22
rect 220 -30 224 -22
rect -55 -34 -48 -30
rect -44 -34 -27 -30
rect -23 -34 -11 -30
rect -7 -34 4 -30
rect 8 -34 29 -30
rect 33 -34 50 -30
rect 54 -34 66 -30
rect 70 -34 81 -30
rect 85 -34 106 -30
rect 110 -34 127 -30
rect 131 -34 143 -30
rect 147 -34 158 -30
rect 162 -34 183 -30
rect 187 -34 204 -30
rect 208 -34 220 -30
rect 224 -34 235 -30
rect 239 -34 242 -30
<< ntransistor >>
rect -45 -24 -42 -16
rect -30 -24 -27 -16
rect -3 -24 -1 -16
rect 32 -24 35 -16
rect 47 -24 50 -16
rect 74 -24 76 -16
rect 109 -24 112 -16
rect 124 -24 127 -16
rect 151 -24 153 -16
rect 186 -24 189 -16
rect 201 -24 204 -16
rect 228 -24 230 -16
<< ptransistor >>
rect -45 16 -42 24
rect -30 16 -27 24
rect -3 16 -1 24
rect 32 16 35 24
rect 47 16 50 24
rect 74 16 76 24
rect 109 16 112 24
rect 124 16 127 24
rect 151 16 153 24
rect 186 16 189 24
rect 201 16 204 24
rect 228 16 230 24
<< polycontact >>
rect -7 -3 -3 1
rect 9 -1 13 3
rect 70 -3 74 1
rect 86 -1 90 3
rect 147 -3 151 1
rect 163 -1 167 3
rect 224 -3 228 1
rect 240 -1 244 3
<< ndcontact >>
rect -53 -22 -49 -18
rect -23 -22 -19 -18
rect -11 -22 -7 -18
rect 3 -22 7 -18
rect 24 -22 28 -18
rect 54 -22 58 -18
rect 66 -22 70 -18
rect 80 -22 84 -18
rect 101 -22 105 -18
rect 131 -22 135 -18
rect 143 -22 147 -18
rect 157 -22 161 -18
rect 178 -22 182 -18
rect 208 -22 212 -18
rect 220 -22 224 -18
rect 234 -22 238 -18
<< pdcontact >>
rect -53 18 -49 22
rect -38 18 -34 22
rect -23 18 -19 22
rect -11 18 -7 22
rect 3 18 7 22
rect 24 18 28 22
rect 39 18 43 22
rect 54 18 58 22
rect 66 18 70 22
rect 80 18 84 22
rect 101 18 105 22
rect 116 18 120 22
rect 131 18 135 22
rect 143 18 147 22
rect 157 18 161 22
rect 178 18 182 22
rect 193 18 197 22
rect 208 18 212 22
rect 220 18 224 22
rect 234 18 238 22
<< nbccdiffcontact >>
rect -11 32 -7 36
rect 66 32 70 36
rect 143 32 147 36
rect 220 32 224 36
<< psubstratepcontact >>
rect -48 -34 -44 -30
rect -27 -34 -23 -30
rect -11 -34 -7 -30
rect 4 -34 8 -30
rect 29 -34 33 -30
rect 50 -34 54 -30
rect 66 -34 70 -30
rect 81 -34 85 -30
rect 106 -34 110 -30
rect 127 -34 131 -30
rect 143 -34 147 -30
rect 158 -34 162 -30
rect 183 -34 187 -30
rect 204 -34 208 -30
rect 220 -34 224 -30
rect 235 -34 239 -30
<< nsubstratencontact >>
rect -48 32 -44 36
rect -29 32 -25 36
rect 3 32 7 36
rect 29 32 33 36
rect 48 32 52 36
rect 80 32 84 36
rect 106 32 110 36
rect 125 32 129 36
rect 157 32 161 36
rect 183 32 187 36
rect 202 32 206 36
rect 234 32 238 36
<< labels >>
rlabel polysilicon -40 56 -40 56 5 a0
rlabel polysilicon -31 56 -31 56 5 b0
rlabel polysilicon 37 55 37 55 5 a1
rlabel polysilicon 46 55 46 55 5 b1
rlabel polysilicon 114 55 114 55 5 a2
rlabel polysilicon 123 55 123 55 5 b2
rlabel polysilicon 191 55 191 55 5 a3
rlabel polysilicon 200 55 200 55 5 b3
rlabel polysilicon 13 -46 13 -46 1 s0
rlabel polysilicon 90 -46 90 -46 1 s1
rlabel polysilicon 167 -46 167 -46 1 s2
rlabel polysilicon 244 -46 244 -46 8 s3
rlabel metal1 98 -32 98 -32 1 gnd
rlabel metal1 99 34 99 34 1 Vdd
<< end >>
