magic
tech scmos
timestamp 1700586729
<< nwell >>
rect -66 49 61 61
<< polysilicon >>
rect -54 59 -51 63
rect -30 59 -27 63
rect -4 59 -1 63
rect 20 59 23 63
rect 47 59 49 63
rect -54 18 -51 51
rect -30 18 -27 51
rect -4 18 -1 51
rect 20 18 23 51
rect 47 18 49 51
rect -54 8 -51 10
rect -30 8 -27 10
rect -4 8 -1 10
rect 20 8 23 10
rect 47 8 49 10
<< ndiffusion >>
rect -64 16 -54 18
rect -64 12 -62 16
rect -58 12 -54 16
rect -64 10 -54 12
rect -51 16 -44 18
rect -51 12 -48 16
rect -51 10 -44 12
rect -40 16 -30 18
rect -40 12 -38 16
rect -34 12 -30 16
rect -40 10 -30 12
rect -27 16 -18 18
rect -27 12 -24 16
rect -20 12 -18 16
rect -27 10 -18 12
rect -14 16 -4 18
rect -14 12 -12 16
rect -8 12 -4 16
rect -14 10 -4 12
rect -1 16 7 18
rect -1 12 2 16
rect 6 12 7 16
rect -1 10 7 12
rect 11 16 20 18
rect 11 12 12 16
rect 16 12 20 16
rect 11 10 20 12
rect 23 16 33 18
rect 23 12 27 16
rect 31 12 33 16
rect 23 10 33 12
rect 37 16 47 18
rect 37 12 39 16
rect 43 12 47 16
rect 37 10 47 12
rect 49 16 59 18
rect 49 12 53 16
rect 57 12 59 16
rect 49 10 59 12
<< pdiffusion >>
rect -64 57 -54 59
rect -64 53 -62 57
rect -58 53 -54 57
rect -64 51 -54 53
rect -51 51 -30 59
rect -27 51 -4 59
rect -1 51 20 59
rect 23 57 33 59
rect 23 53 27 57
rect 31 53 33 57
rect 23 51 33 53
rect 37 57 47 59
rect 37 53 39 57
rect 43 53 47 57
rect 37 51 47 53
rect 49 57 59 59
rect 49 53 53 57
rect 57 53 59 57
rect 49 51 59 53
<< metal1 >>
rect -66 67 -57 71
rect -53 67 -33 71
rect -29 67 -7 71
rect -3 67 21 71
rect 25 67 39 71
rect 43 67 53 71
rect 57 67 61 71
rect -62 57 -58 67
rect 39 57 43 67
rect -66 42 16 46
rect -66 35 -8 39
rect 27 36 31 53
rect 53 38 57 53
rect 2 32 43 36
rect 53 34 61 38
rect -66 28 -34 32
rect 2 25 6 32
rect -66 21 -58 25
rect -48 21 6 25
rect -48 16 -44 21
rect -24 16 -20 21
rect 2 16 6 21
rect 27 16 31 32
rect 53 16 57 34
rect -62 4 -58 12
rect -38 4 -34 12
rect -12 4 -8 12
rect 12 4 16 12
rect 39 4 43 12
rect -64 0 -57 4
rect -53 0 -33 4
rect -29 0 -7 4
rect -3 0 23 4
rect 27 0 39 4
rect 43 0 54 4
rect 58 0 61 4
<< ntransistor >>
rect -54 10 -51 18
rect -30 10 -27 18
rect -4 10 -1 18
rect 20 10 23 18
rect 47 10 49 18
<< ptransistor >>
rect -54 51 -51 59
rect -30 51 -27 59
rect -4 51 -1 59
rect 20 51 23 59
rect 47 51 49 59
<< polycontact >>
rect -58 21 -54 25
rect -34 28 -30 32
rect -8 35 -4 39
rect 16 42 20 46
rect 43 32 47 36
<< ndcontact >>
rect -62 12 -58 16
rect -48 12 -44 16
rect -38 12 -34 16
rect -24 12 -20 16
rect -12 12 -8 16
rect 2 12 6 16
rect 12 12 16 16
rect 27 12 31 16
rect 39 12 43 16
rect 53 12 57 16
<< pdcontact >>
rect -62 53 -58 57
rect 27 53 31 57
rect 39 53 43 57
rect 53 53 57 57
<< nbccdiffcontact >>
rect 39 67 43 71
<< psubstratepcontact >>
rect -57 0 -53 4
rect -33 0 -29 4
rect -7 0 -3 4
rect 23 0 27 4
rect 39 0 43 4
rect 54 0 58 4
<< nsubstratencontact >>
rect -57 67 -53 71
rect -33 67 -29 71
rect -7 67 -3 71
rect 21 67 25 71
rect 53 67 57 71
<< end >>
