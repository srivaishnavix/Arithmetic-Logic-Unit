* SPICE3 file created from 3ANDGAT.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'


.option scale=1u

M1000 a_31_52# Va Vdd w_16_50# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1001 Vout a_31_52# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1002 Vout a_31_52# Vdd w_16_50# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1003 a_46_11# Vb a_31_11# Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=48p ps=20u
M1004 a_31_52# Vc a_46_11# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1005 a_31_52# Vb a_31_52# w_16_50# CMOSP w=8 l=3
+  ad=48p pd=20u as=0.192n ps=80u
M1006 Vdd Vc a_31_52# w_16_50# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1007 a_31_11# Va gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
C0 gnd 0 14.476f 
C1 Vout 0 6.58f 
C2 a_31_52# 0 24.354f 
C3 Vc 0 19.431f 
C4 Vb 0 17.175001f 
C5 Va 0 14.919f 
C6 Vdd 0 15.98f 


Va Va gnd 1
Vb Vb gnd 1
Vc Vc gnd 0



.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(Va) v(Vb)+2 v(Vc)+4 v(Vout)+6
.end
.endc