magic
tech scmos
timestamp 1701025380
<< nwell >>
rect 1390 297 1517 309
rect 757 198 851 210
rect 864 198 947 210
rect 1089 206 1183 218
rect 1192 206 1290 218
rect 412 185 506 197
rect 515 185 583 197
rect 66 142 160 154
rect 1471 133 1569 145
rect 96 47 138 59
rect 442 50 484 62
rect 800 55 842 67
rect 1144 63 1186 75
rect 29 8 71 20
rect 164 12 206 24
rect 237 3 263 15
rect 375 11 417 23
rect 510 15 552 27
rect 583 6 609 18
rect 733 16 775 28
rect 868 20 910 32
rect 1077 24 1119 36
rect 1212 28 1254 40
rect 941 11 967 23
rect 1285 19 1311 31
rect 96 -36 138 -24
rect 442 -33 484 -21
rect 800 -28 842 -16
rect 1144 -20 1186 -8
rect 74 -138 168 -126
rect 729 -167 823 -155
rect 836 -167 919 -155
rect 1075 -165 1169 -153
rect 1178 -165 1276 -153
rect 404 -182 498 -170
rect 507 -182 574 -170
rect 1337 -366 1464 -354
<< polysilicon >>
rect 1402 307 1405 311
rect 1426 307 1429 311
rect 1452 307 1455 311
rect 1476 307 1479 311
rect 1503 307 1505 311
rect 179 290 1337 294
rect 597 283 1335 287
rect 966 276 1333 280
rect 1402 266 1405 299
rect 1426 266 1429 299
rect 1452 266 1455 299
rect 1476 266 1479 299
rect 1503 266 1505 299
rect 1402 256 1405 258
rect 1426 256 1429 258
rect 1452 256 1455 258
rect 1476 256 1479 258
rect 1503 256 1505 258
rect 1101 216 1103 220
rect 1127 216 1130 220
rect 1142 216 1145 220
rect 1169 216 1171 220
rect 1204 216 1207 220
rect 1219 216 1222 220
rect 1234 216 1237 220
rect 1249 216 1252 220
rect 1276 216 1278 220
rect 769 208 771 212
rect 795 208 798 212
rect 810 208 813 212
rect 837 208 839 212
rect 876 208 879 212
rect 891 208 894 212
rect 906 208 909 212
rect 933 208 935 212
rect 424 195 426 199
rect 450 195 453 199
rect 465 195 468 199
rect 492 195 494 199
rect 527 195 530 199
rect 542 195 545 199
rect 569 195 571 199
rect 680 189 755 193
rect 322 176 410 180
rect 339 159 410 163
rect 78 152 80 156
rect 104 152 107 156
rect 119 152 122 156
rect 146 152 148 156
rect 424 155 426 187
rect 450 164 453 187
rect 465 172 468 187
rect 464 168 468 172
rect 449 160 453 164
rect 450 155 453 160
rect 465 155 468 168
rect 492 155 494 187
rect 527 164 530 187
rect 542 172 545 187
rect 541 168 545 172
rect 509 160 530 164
rect 424 145 426 147
rect 450 145 453 147
rect 465 145 468 147
rect 492 145 494 147
rect -24 133 64 137
rect -7 116 64 120
rect 78 112 80 144
rect 104 121 107 144
rect 119 129 122 144
rect 118 125 122 129
rect 103 117 107 121
rect 104 112 107 117
rect 119 112 122 125
rect 146 112 148 144
rect 509 134 513 160
rect 527 155 530 160
rect 542 155 545 168
rect 569 155 571 187
rect 697 172 755 176
rect 769 168 771 200
rect 795 177 798 200
rect 810 185 813 200
rect 809 181 813 185
rect 794 173 798 177
rect 795 168 798 173
rect 810 168 813 181
rect 837 168 839 200
rect 876 167 879 200
rect 891 167 894 200
rect 906 167 909 200
rect 933 167 935 200
rect 1024 197 1087 201
rect 1041 180 1087 184
rect 1101 176 1103 208
rect 1127 185 1130 208
rect 1142 193 1145 208
rect 1141 189 1145 193
rect 1126 181 1130 185
rect 1127 176 1130 181
rect 1142 176 1145 189
rect 1169 176 1171 208
rect 1204 175 1207 208
rect 1219 175 1222 208
rect 1234 175 1237 208
rect 1249 175 1252 208
rect 1276 175 1278 208
rect 769 158 771 160
rect 795 158 798 160
rect 810 158 813 160
rect 837 158 839 160
rect 1101 166 1103 168
rect 1127 166 1130 168
rect 1142 166 1145 168
rect 1169 166 1171 168
rect 1204 165 1207 167
rect 876 157 879 159
rect 527 145 530 147
rect 542 145 545 147
rect 569 145 571 147
rect 891 134 894 159
rect 906 158 909 159
rect 902 155 909 158
rect 933 157 935 159
rect 902 146 905 155
rect 1219 134 1222 167
rect 1234 144 1237 167
rect 1249 165 1252 167
rect 1276 165 1278 167
rect 1244 162 1252 165
rect 1244 144 1247 162
rect 1483 143 1486 147
rect 1498 143 1501 147
rect 1513 143 1516 147
rect 1528 143 1531 147
rect 1555 143 1557 147
rect 292 130 1440 134
rect 1436 126 1467 130
rect 639 122 902 124
rect 906 122 1234 124
rect 1238 123 1441 124
rect 1238 122 1467 123
rect 639 120 1467 122
rect 1436 119 1467 120
rect 985 113 1244 115
rect 1436 115 1467 116
rect 1248 113 1467 115
rect 985 112 1467 113
rect 985 111 1442 112
rect 1443 105 1467 109
rect 78 102 80 104
rect 104 102 107 104
rect 119 102 122 104
rect 146 102 148 104
rect 1443 101 1447 105
rect 1483 102 1486 135
rect 1498 102 1501 135
rect 1513 102 1516 135
rect 1528 102 1531 135
rect 1555 102 1557 135
rect 1333 97 1447 101
rect 1156 73 1159 77
rect 1171 73 1174 77
rect 812 65 815 69
rect 827 65 830 69
rect 108 57 111 61
rect 123 57 126 61
rect 454 60 457 64
rect 469 60 472 64
rect 108 26 111 49
rect 123 34 126 49
rect 122 30 126 34
rect 107 22 111 26
rect 41 18 44 22
rect 56 18 59 22
rect 108 17 111 22
rect 123 17 126 30
rect 454 29 457 52
rect 469 37 472 52
rect 468 33 472 37
rect 812 34 815 57
rect 827 42 830 57
rect 1156 42 1159 65
rect 1171 50 1174 65
rect 1170 46 1174 50
rect 826 38 830 42
rect 1155 38 1159 42
rect 176 22 179 26
rect 191 22 194 26
rect 453 25 457 29
rect -24 -9 8 -5
rect 41 -13 44 10
rect 56 -5 59 10
rect 387 21 390 25
rect 402 21 405 25
rect 108 7 111 9
rect 123 7 126 9
rect 55 -9 59 -5
rect 176 -9 179 14
rect 191 -1 194 14
rect 249 13 251 17
rect 454 20 457 25
rect 469 20 472 33
rect 811 30 815 34
rect 522 25 525 29
rect 537 25 540 29
rect 190 -5 194 -1
rect -7 -17 8 -13
rect 40 -17 44 -13
rect 41 -22 44 -17
rect 56 -22 59 -9
rect 175 -13 179 -9
rect 176 -18 179 -13
rect 191 -18 194 -5
rect 249 -9 251 5
rect 322 -6 354 -2
rect 387 -10 390 13
rect 402 -2 405 13
rect 745 26 748 30
rect 760 26 763 30
rect 454 10 457 12
rect 469 10 472 12
rect 401 -6 405 -2
rect 522 -6 525 17
rect 537 2 540 17
rect 595 16 597 20
rect 812 25 815 30
rect 827 25 830 38
rect 1089 34 1092 38
rect 1104 34 1107 38
rect 880 30 883 34
rect 895 30 898 34
rect 536 -2 540 2
rect 339 -14 354 -10
rect 386 -14 390 -10
rect 108 -26 111 -22
rect 123 -26 126 -22
rect 249 -19 251 -17
rect 387 -19 390 -14
rect 402 -19 405 -6
rect 521 -10 525 -6
rect 522 -15 525 -10
rect 537 -15 540 -2
rect 595 -6 597 8
rect 680 -1 712 3
rect 745 -5 748 18
rect 760 3 763 18
rect 1156 33 1159 38
rect 1171 33 1174 46
rect 1224 38 1227 42
rect 1239 38 1242 42
rect 812 15 815 17
rect 827 15 830 17
rect 759 -1 763 3
rect 880 -1 883 22
rect 895 7 898 22
rect 953 21 955 25
rect 894 3 898 7
rect 697 -9 712 -5
rect 744 -9 748 -5
rect 745 -14 748 -9
rect 760 -14 763 -1
rect 879 -5 883 -1
rect 880 -10 883 -5
rect 895 -10 898 3
rect 953 -1 955 13
rect 1024 7 1056 11
rect 1089 3 1092 26
rect 1104 11 1107 26
rect 1156 23 1159 25
rect 1171 23 1174 25
rect 1103 7 1107 11
rect 1224 7 1227 30
rect 1239 15 1242 30
rect 1297 29 1299 33
rect 1238 11 1242 15
rect 1041 -1 1056 3
rect 1088 -1 1092 3
rect 1089 -6 1092 -1
rect 1104 -6 1107 7
rect 1223 3 1227 7
rect 1224 -2 1227 3
rect 1239 -2 1242 11
rect 1297 7 1299 21
rect 1333 16 1337 97
rect 1483 92 1486 94
rect 1498 92 1501 94
rect 1513 92 1516 94
rect 1528 92 1531 94
rect 1555 92 1557 94
rect 1317 12 1337 16
rect 41 -32 44 -30
rect 56 -32 59 -30
rect 176 -28 179 -26
rect 191 -28 194 -26
rect 454 -23 457 -19
rect 469 -23 472 -19
rect 595 -16 597 -14
rect 387 -29 390 -27
rect 402 -29 405 -27
rect 522 -25 525 -23
rect 537 -25 540 -23
rect 812 -18 815 -14
rect 827 -18 830 -14
rect 953 -11 955 -9
rect 1156 -10 1159 -6
rect 1171 -10 1174 -6
rect 1297 -3 1299 -1
rect 745 -24 748 -22
rect 760 -24 763 -22
rect 880 -20 883 -18
rect 895 -20 898 -18
rect 1089 -16 1092 -14
rect 1104 -16 1107 -14
rect 1224 -12 1227 -10
rect 1239 -12 1242 -10
rect 108 -57 111 -34
rect 123 -49 126 -34
rect 122 -53 126 -49
rect 107 -61 111 -57
rect 108 -66 111 -61
rect 123 -66 126 -53
rect 454 -54 457 -31
rect 469 -46 472 -31
rect 468 -50 472 -46
rect 812 -49 815 -26
rect 827 -41 830 -26
rect 1156 -41 1159 -18
rect 1171 -33 1174 -18
rect 1170 -37 1174 -33
rect 826 -45 830 -41
rect 1155 -45 1159 -41
rect 453 -58 457 -54
rect 454 -63 457 -58
rect 469 -63 472 -50
rect 811 -53 815 -49
rect 812 -58 815 -53
rect 827 -58 830 -45
rect 1156 -50 1159 -45
rect 1171 -50 1174 -37
rect 1156 -60 1159 -58
rect 1171 -60 1174 -58
rect 812 -68 815 -66
rect 827 -68 830 -66
rect 454 -73 457 -71
rect 469 -73 472 -71
rect 108 -76 111 -74
rect 123 -76 126 -74
rect 86 -128 88 -124
rect 112 -128 115 -124
rect 127 -128 130 -124
rect 154 -128 156 -124
rect -7 -147 72 -143
rect -24 -164 72 -160
rect 86 -168 88 -136
rect 112 -159 115 -136
rect 127 -151 130 -136
rect 126 -155 130 -151
rect 111 -163 115 -159
rect 112 -168 115 -163
rect 127 -168 130 -155
rect 154 -168 156 -136
rect 741 -157 743 -153
rect 767 -157 770 -153
rect 782 -157 785 -153
rect 809 -157 811 -153
rect 848 -157 851 -153
rect 863 -157 866 -153
rect 878 -157 881 -153
rect 905 -157 907 -153
rect 1087 -155 1089 -151
rect 1113 -155 1116 -151
rect 1128 -155 1131 -151
rect 1155 -155 1157 -151
rect 1190 -155 1193 -151
rect 1205 -155 1208 -151
rect 1220 -155 1223 -151
rect 1235 -155 1238 -151
rect 1262 -155 1264 -151
rect 416 -172 418 -168
rect 442 -172 445 -168
rect 457 -172 460 -168
rect 484 -172 486 -168
rect 519 -172 522 -168
rect 534 -172 537 -168
rect 561 -172 563 -168
rect 86 -178 88 -176
rect 112 -178 115 -176
rect 127 -178 130 -176
rect 154 -178 156 -176
rect 697 -176 727 -172
rect 339 -191 402 -187
rect 322 -208 402 -204
rect 416 -212 418 -180
rect 442 -203 445 -180
rect 457 -195 460 -180
rect 456 -199 460 -195
rect 441 -207 445 -203
rect 442 -212 445 -207
rect 457 -212 460 -199
rect 484 -212 486 -180
rect 519 -203 522 -180
rect 534 -195 537 -180
rect 533 -199 537 -195
rect 501 -207 522 -203
rect 416 -222 418 -220
rect 442 -222 445 -220
rect 457 -222 460 -220
rect 484 -222 486 -220
rect 501 -275 505 -207
rect 519 -212 522 -207
rect 534 -212 537 -199
rect 561 -212 563 -180
rect 680 -193 727 -189
rect 741 -197 743 -165
rect 767 -188 770 -165
rect 782 -180 785 -165
rect 781 -184 785 -180
rect 766 -192 770 -188
rect 767 -197 770 -192
rect 782 -197 785 -184
rect 809 -197 811 -165
rect 848 -198 851 -165
rect 863 -198 866 -165
rect 878 -198 881 -165
rect 905 -198 907 -165
rect 1041 -174 1073 -170
rect 1024 -191 1073 -187
rect 1087 -195 1089 -163
rect 1113 -186 1116 -163
rect 1128 -178 1131 -163
rect 1127 -182 1131 -178
rect 1112 -190 1116 -186
rect 1113 -195 1116 -190
rect 1128 -195 1131 -182
rect 1155 -195 1157 -163
rect 741 -207 743 -205
rect 767 -207 770 -205
rect 782 -207 785 -205
rect 809 -207 811 -205
rect 1190 -196 1193 -163
rect 1205 -196 1208 -163
rect 1220 -196 1223 -163
rect 1235 -196 1238 -163
rect 1262 -196 1264 -163
rect 1087 -205 1089 -203
rect 1113 -205 1116 -203
rect 1128 -205 1131 -203
rect 1155 -205 1157 -203
rect 1190 -206 1193 -204
rect 848 -208 851 -206
rect 519 -222 522 -220
rect 534 -222 537 -220
rect 561 -222 563 -220
rect 863 -266 866 -206
rect 878 -207 881 -206
rect 874 -210 881 -207
rect 905 -208 907 -206
rect 874 -220 877 -210
rect 874 -223 881 -220
rect 878 -251 881 -223
rect 878 -253 882 -251
rect 1205 -256 1208 -204
rect 1220 -243 1223 -204
rect 1235 -206 1238 -204
rect 1262 -206 1264 -204
rect 1230 -209 1238 -206
rect 1230 -215 1233 -209
rect 1230 -218 1238 -215
rect 1235 -243 1238 -218
rect 985 -260 1331 -256
rect 639 -268 1220 -266
rect 1224 -268 1331 -266
rect 639 -270 1331 -268
rect 296 -277 878 -275
rect 882 -277 1235 -275
rect 1239 -277 1334 -275
rect 296 -279 1334 -277
rect 1349 -356 1352 -352
rect 1373 -356 1376 -352
rect 1399 -356 1402 -352
rect 1423 -356 1426 -352
rect 1450 -356 1452 -352
rect 1349 -397 1352 -364
rect 1373 -397 1376 -364
rect 1399 -397 1402 -364
rect 1423 -397 1426 -364
rect 1450 -397 1452 -364
rect 1349 -407 1352 -405
rect 1373 -407 1376 -405
rect 1399 -407 1402 -405
rect 1423 -407 1426 -405
rect 1450 -407 1452 -405
<< ndiffusion >>
rect 1392 264 1402 266
rect 1392 260 1394 264
rect 1398 260 1402 264
rect 1392 258 1402 260
rect 1405 264 1412 266
rect 1405 260 1408 264
rect 1405 258 1412 260
rect 1416 264 1426 266
rect 1416 260 1418 264
rect 1422 260 1426 264
rect 1416 258 1426 260
rect 1429 264 1438 266
rect 1429 260 1432 264
rect 1436 260 1438 264
rect 1429 258 1438 260
rect 1442 264 1452 266
rect 1442 260 1444 264
rect 1448 260 1452 264
rect 1442 258 1452 260
rect 1455 264 1463 266
rect 1455 260 1458 264
rect 1462 260 1463 264
rect 1455 258 1463 260
rect 1467 264 1476 266
rect 1467 260 1468 264
rect 1472 260 1476 264
rect 1467 258 1476 260
rect 1479 264 1489 266
rect 1479 260 1483 264
rect 1487 260 1489 264
rect 1479 258 1489 260
rect 1493 264 1503 266
rect 1493 260 1495 264
rect 1499 260 1503 264
rect 1493 258 1503 260
rect 1505 264 1515 266
rect 1505 260 1509 264
rect 1513 260 1515 264
rect 1505 258 1515 260
rect 414 153 424 155
rect 414 149 416 153
rect 420 149 424 153
rect 414 147 424 149
rect 426 153 436 155
rect 426 149 430 153
rect 434 149 436 153
rect 426 147 436 149
rect 440 153 450 155
rect 440 149 442 153
rect 446 149 450 153
rect 440 147 450 149
rect 453 147 465 155
rect 468 153 478 155
rect 468 149 472 153
rect 476 149 478 153
rect 468 147 478 149
rect 482 153 492 155
rect 482 149 484 153
rect 488 149 492 153
rect 482 147 492 149
rect 494 153 504 155
rect 494 149 498 153
rect 502 149 504 153
rect 494 147 504 149
rect 759 166 769 168
rect 759 162 761 166
rect 765 162 769 166
rect 759 160 769 162
rect 771 166 781 168
rect 771 162 775 166
rect 779 162 781 166
rect 771 160 781 162
rect 785 166 795 168
rect 785 162 787 166
rect 791 162 795 166
rect 785 160 795 162
rect 798 160 810 168
rect 813 166 823 168
rect 813 162 817 166
rect 821 162 823 166
rect 813 160 823 162
rect 827 166 837 168
rect 827 162 829 166
rect 833 162 837 166
rect 827 160 837 162
rect 839 166 849 168
rect 1091 174 1101 176
rect 1091 170 1093 174
rect 1097 170 1101 174
rect 1091 168 1101 170
rect 1103 174 1113 176
rect 1103 170 1107 174
rect 1111 170 1113 174
rect 1103 168 1113 170
rect 1117 174 1127 176
rect 1117 170 1119 174
rect 1123 170 1127 174
rect 1117 168 1127 170
rect 1130 168 1142 176
rect 1145 174 1155 176
rect 1145 170 1149 174
rect 1153 170 1155 174
rect 1145 168 1155 170
rect 1159 174 1169 176
rect 1159 170 1161 174
rect 1165 170 1169 174
rect 1159 168 1169 170
rect 1171 174 1181 176
rect 1171 170 1175 174
rect 1179 170 1181 174
rect 1171 168 1181 170
rect 1194 173 1204 175
rect 1194 169 1196 173
rect 1200 169 1204 173
rect 839 162 843 166
rect 847 162 849 166
rect 839 160 849 162
rect 866 165 876 167
rect 866 161 868 165
rect 872 161 876 165
rect 866 159 876 161
rect 879 159 891 167
rect 894 159 906 167
rect 909 165 919 167
rect 909 161 913 165
rect 917 161 919 165
rect 909 159 919 161
rect 923 165 933 167
rect 923 161 925 165
rect 929 161 933 165
rect 923 159 933 161
rect 935 165 945 167
rect 1194 167 1204 169
rect 1207 167 1219 175
rect 1222 167 1234 175
rect 1237 167 1249 175
rect 1252 173 1262 175
rect 1252 169 1256 173
rect 1260 169 1262 173
rect 1252 167 1262 169
rect 1266 173 1276 175
rect 1266 169 1268 173
rect 1272 169 1276 173
rect 1266 167 1276 169
rect 1278 173 1288 175
rect 1278 169 1282 173
rect 1286 169 1288 173
rect 1278 167 1288 169
rect 935 161 939 165
rect 943 161 945 165
rect 935 159 945 161
rect 517 153 527 155
rect 517 149 519 153
rect 523 149 527 153
rect 517 147 527 149
rect 530 147 542 155
rect 545 153 555 155
rect 545 149 549 153
rect 553 149 555 153
rect 545 147 555 149
rect 559 153 569 155
rect 559 149 561 153
rect 565 149 569 153
rect 559 147 569 149
rect 571 153 581 155
rect 571 149 575 153
rect 579 149 581 153
rect 571 147 581 149
rect 68 110 78 112
rect 68 106 70 110
rect 74 106 78 110
rect 68 104 78 106
rect 80 110 90 112
rect 80 106 84 110
rect 88 106 90 110
rect 80 104 90 106
rect 94 110 104 112
rect 94 106 96 110
rect 100 106 104 110
rect 94 104 104 106
rect 107 104 119 112
rect 122 110 132 112
rect 122 106 126 110
rect 130 106 132 110
rect 122 104 132 106
rect 136 110 146 112
rect 136 106 138 110
rect 142 106 146 110
rect 136 104 146 106
rect 148 110 158 112
rect 148 106 152 110
rect 156 106 158 110
rect 148 104 158 106
rect 1473 100 1483 102
rect 98 15 108 17
rect 98 11 100 15
rect 104 11 108 15
rect 98 9 108 11
rect 111 9 123 17
rect 126 15 136 17
rect 126 11 130 15
rect 134 11 136 15
rect 126 9 136 11
rect 444 18 454 20
rect 444 14 446 18
rect 450 14 454 18
rect 239 -11 249 -9
rect 239 -15 241 -11
rect 245 -15 249 -11
rect 239 -17 249 -15
rect 251 -11 261 -9
rect 444 12 454 14
rect 457 12 469 20
rect 472 18 482 20
rect 472 14 476 18
rect 480 14 482 18
rect 472 12 482 14
rect 802 23 812 25
rect 802 19 804 23
rect 808 19 812 23
rect 251 -15 255 -11
rect 259 -15 261 -11
rect 251 -17 261 -15
rect 166 -20 176 -18
rect 31 -24 41 -22
rect 31 -28 33 -24
rect 37 -28 41 -24
rect 31 -30 41 -28
rect 44 -30 56 -22
rect 59 -24 69 -22
rect 59 -28 63 -24
rect 67 -28 69 -24
rect 166 -24 168 -20
rect 172 -24 176 -20
rect 166 -26 176 -24
rect 179 -26 191 -18
rect 194 -20 204 -18
rect 802 17 812 19
rect 815 17 827 25
rect 830 23 840 25
rect 830 19 834 23
rect 838 19 840 23
rect 1146 31 1156 33
rect 1146 27 1148 31
rect 1152 27 1156 31
rect 830 17 840 19
rect 585 -8 595 -6
rect 585 -12 587 -8
rect 591 -12 595 -8
rect 585 -14 595 -12
rect 597 -8 607 -6
rect 597 -12 601 -8
rect 605 -12 607 -8
rect 597 -14 607 -12
rect 1146 25 1156 27
rect 1159 25 1171 33
rect 1174 31 1184 33
rect 1174 27 1178 31
rect 1182 27 1184 31
rect 1174 25 1184 27
rect 943 -3 953 -1
rect 943 -7 945 -3
rect 949 -7 953 -3
rect 943 -9 953 -7
rect 955 -3 965 -1
rect 955 -7 959 -3
rect 963 -7 965 -3
rect 1473 96 1475 100
rect 1479 96 1483 100
rect 1473 94 1483 96
rect 1486 94 1498 102
rect 1501 94 1513 102
rect 1516 94 1528 102
rect 1531 100 1541 102
rect 1531 96 1535 100
rect 1539 96 1541 100
rect 1531 94 1541 96
rect 1545 100 1555 102
rect 1545 96 1547 100
rect 1551 96 1555 100
rect 1545 94 1555 96
rect 1557 100 1567 102
rect 1557 96 1561 100
rect 1565 96 1567 100
rect 1557 94 1567 96
rect 1287 5 1297 7
rect 1287 1 1289 5
rect 1293 1 1297 5
rect 1287 -1 1297 1
rect 1299 5 1309 7
rect 1299 1 1303 5
rect 1307 1 1309 5
rect 1299 -1 1309 1
rect 1214 -4 1224 -2
rect 955 -9 965 -7
rect 1079 -8 1089 -6
rect 870 -12 880 -10
rect 512 -17 522 -15
rect 194 -24 198 -20
rect 202 -24 204 -20
rect 377 -21 387 -19
rect 194 -26 204 -24
rect 59 -30 69 -28
rect 377 -25 379 -21
rect 383 -25 387 -21
rect 377 -27 387 -25
rect 390 -27 402 -19
rect 405 -21 415 -19
rect 405 -25 409 -21
rect 413 -25 415 -21
rect 512 -21 514 -17
rect 518 -21 522 -17
rect 512 -23 522 -21
rect 525 -23 537 -15
rect 540 -17 550 -15
rect 735 -16 745 -14
rect 540 -21 544 -17
rect 548 -21 550 -17
rect 735 -20 737 -16
rect 741 -20 745 -16
rect 540 -23 550 -21
rect 405 -27 415 -25
rect 735 -22 745 -20
rect 748 -22 760 -14
rect 763 -16 773 -14
rect 763 -20 767 -16
rect 771 -20 773 -16
rect 870 -16 872 -12
rect 876 -16 880 -12
rect 870 -18 880 -16
rect 883 -18 895 -10
rect 898 -12 908 -10
rect 898 -16 902 -12
rect 906 -16 908 -12
rect 1079 -12 1081 -8
rect 1085 -12 1089 -8
rect 1079 -14 1089 -12
rect 1092 -14 1104 -6
rect 1107 -8 1117 -6
rect 1107 -12 1111 -8
rect 1115 -12 1117 -8
rect 1214 -8 1216 -4
rect 1220 -8 1224 -4
rect 1214 -10 1224 -8
rect 1227 -10 1239 -2
rect 1242 -4 1252 -2
rect 1242 -8 1246 -4
rect 1250 -8 1252 -4
rect 1242 -10 1252 -8
rect 1107 -14 1117 -12
rect 898 -18 908 -16
rect 763 -22 773 -20
rect 1146 -52 1156 -50
rect 1146 -56 1148 -52
rect 1152 -56 1156 -52
rect 1146 -58 1156 -56
rect 1159 -58 1171 -50
rect 1174 -52 1184 -50
rect 1174 -56 1178 -52
rect 1182 -56 1184 -52
rect 1174 -58 1184 -56
rect 802 -60 812 -58
rect 444 -65 454 -63
rect 98 -68 108 -66
rect 98 -72 100 -68
rect 104 -72 108 -68
rect 98 -74 108 -72
rect 111 -74 123 -66
rect 126 -68 136 -66
rect 126 -72 130 -68
rect 134 -72 136 -68
rect 444 -69 446 -65
rect 450 -69 454 -65
rect 444 -71 454 -69
rect 457 -71 469 -63
rect 472 -65 482 -63
rect 472 -69 476 -65
rect 480 -69 482 -65
rect 802 -64 804 -60
rect 808 -64 812 -60
rect 802 -66 812 -64
rect 815 -66 827 -58
rect 830 -60 840 -58
rect 830 -64 834 -60
rect 838 -64 840 -60
rect 830 -66 840 -64
rect 472 -71 482 -69
rect 126 -74 136 -72
rect 76 -170 86 -168
rect 76 -174 78 -170
rect 82 -174 86 -170
rect 76 -176 86 -174
rect 88 -170 98 -168
rect 88 -174 92 -170
rect 96 -174 98 -170
rect 88 -176 98 -174
rect 102 -170 112 -168
rect 102 -174 104 -170
rect 108 -174 112 -170
rect 102 -176 112 -174
rect 115 -176 127 -168
rect 130 -170 140 -168
rect 130 -174 134 -170
rect 138 -174 140 -170
rect 130 -176 140 -174
rect 144 -170 154 -168
rect 144 -174 146 -170
rect 150 -174 154 -170
rect 144 -176 154 -174
rect 156 -170 166 -168
rect 156 -174 160 -170
rect 164 -174 166 -170
rect 156 -176 166 -174
rect 406 -214 416 -212
rect 406 -218 408 -214
rect 412 -218 416 -214
rect 406 -220 416 -218
rect 418 -214 428 -212
rect 418 -218 422 -214
rect 426 -218 428 -214
rect 418 -220 428 -218
rect 432 -214 442 -212
rect 432 -218 434 -214
rect 438 -218 442 -214
rect 432 -220 442 -218
rect 445 -220 457 -212
rect 460 -214 470 -212
rect 460 -218 464 -214
rect 468 -218 470 -214
rect 460 -220 470 -218
rect 474 -214 484 -212
rect 474 -218 476 -214
rect 480 -218 484 -214
rect 474 -220 484 -218
rect 486 -214 496 -212
rect 486 -218 490 -214
rect 494 -218 496 -214
rect 486 -220 496 -218
rect 731 -199 741 -197
rect 731 -203 733 -199
rect 737 -203 741 -199
rect 731 -205 741 -203
rect 743 -199 753 -197
rect 743 -203 747 -199
rect 751 -203 753 -199
rect 743 -205 753 -203
rect 757 -199 767 -197
rect 757 -203 759 -199
rect 763 -203 767 -199
rect 757 -205 767 -203
rect 770 -205 782 -197
rect 785 -199 795 -197
rect 785 -203 789 -199
rect 793 -203 795 -199
rect 785 -205 795 -203
rect 799 -199 809 -197
rect 799 -203 801 -199
rect 805 -203 809 -199
rect 799 -205 809 -203
rect 811 -199 821 -197
rect 1077 -197 1087 -195
rect 811 -203 815 -199
rect 819 -203 821 -199
rect 811 -205 821 -203
rect 838 -200 848 -198
rect 838 -204 840 -200
rect 844 -204 848 -200
rect 838 -206 848 -204
rect 851 -206 863 -198
rect 866 -206 878 -198
rect 881 -200 891 -198
rect 881 -204 885 -200
rect 889 -204 891 -200
rect 881 -206 891 -204
rect 895 -200 905 -198
rect 895 -204 897 -200
rect 901 -204 905 -200
rect 895 -206 905 -204
rect 907 -200 917 -198
rect 907 -204 911 -200
rect 915 -204 917 -200
rect 1077 -201 1079 -197
rect 1083 -201 1087 -197
rect 1077 -203 1087 -201
rect 1089 -197 1099 -195
rect 1089 -201 1093 -197
rect 1097 -201 1099 -197
rect 1089 -203 1099 -201
rect 1103 -197 1113 -195
rect 1103 -201 1105 -197
rect 1109 -201 1113 -197
rect 1103 -203 1113 -201
rect 1116 -203 1128 -195
rect 1131 -197 1141 -195
rect 1131 -201 1135 -197
rect 1139 -201 1141 -197
rect 1131 -203 1141 -201
rect 1145 -197 1155 -195
rect 1145 -201 1147 -197
rect 1151 -201 1155 -197
rect 1145 -203 1155 -201
rect 1157 -197 1167 -195
rect 1157 -201 1161 -197
rect 1165 -201 1167 -197
rect 1157 -203 1167 -201
rect 1180 -198 1190 -196
rect 1180 -202 1182 -198
rect 1186 -202 1190 -198
rect 907 -206 917 -204
rect 1180 -204 1190 -202
rect 1193 -204 1205 -196
rect 1208 -204 1220 -196
rect 1223 -204 1235 -196
rect 1238 -198 1248 -196
rect 1238 -202 1242 -198
rect 1246 -202 1248 -198
rect 1238 -204 1248 -202
rect 1252 -198 1262 -196
rect 1252 -202 1254 -198
rect 1258 -202 1262 -198
rect 1252 -204 1262 -202
rect 1264 -198 1274 -196
rect 1264 -202 1268 -198
rect 1272 -202 1274 -198
rect 1264 -204 1274 -202
rect 509 -214 519 -212
rect 509 -218 511 -214
rect 515 -218 519 -214
rect 509 -220 519 -218
rect 522 -220 534 -212
rect 537 -214 547 -212
rect 537 -218 541 -214
rect 545 -218 547 -214
rect 537 -220 547 -218
rect 551 -214 561 -212
rect 551 -218 553 -214
rect 557 -218 561 -214
rect 551 -220 561 -218
rect 563 -214 573 -212
rect 563 -218 567 -214
rect 571 -218 573 -214
rect 563 -220 573 -218
rect 1339 -399 1349 -397
rect 1339 -403 1341 -399
rect 1345 -403 1349 -399
rect 1339 -405 1349 -403
rect 1352 -399 1359 -397
rect 1352 -403 1355 -399
rect 1352 -405 1359 -403
rect 1363 -399 1373 -397
rect 1363 -403 1365 -399
rect 1369 -403 1373 -399
rect 1363 -405 1373 -403
rect 1376 -399 1385 -397
rect 1376 -403 1379 -399
rect 1383 -403 1385 -399
rect 1376 -405 1385 -403
rect 1389 -399 1399 -397
rect 1389 -403 1391 -399
rect 1395 -403 1399 -399
rect 1389 -405 1399 -403
rect 1402 -399 1410 -397
rect 1402 -403 1405 -399
rect 1409 -403 1410 -399
rect 1402 -405 1410 -403
rect 1414 -399 1423 -397
rect 1414 -403 1415 -399
rect 1419 -403 1423 -399
rect 1414 -405 1423 -403
rect 1426 -399 1436 -397
rect 1426 -403 1430 -399
rect 1434 -403 1436 -399
rect 1426 -405 1436 -403
rect 1440 -399 1450 -397
rect 1440 -403 1442 -399
rect 1446 -403 1450 -399
rect 1440 -405 1450 -403
rect 1452 -399 1462 -397
rect 1452 -403 1456 -399
rect 1460 -403 1462 -399
rect 1452 -405 1462 -403
<< pdiffusion >>
rect 1392 305 1402 307
rect 1392 301 1394 305
rect 1398 301 1402 305
rect 1392 299 1402 301
rect 1405 299 1426 307
rect 1429 299 1452 307
rect 1455 299 1476 307
rect 1479 305 1489 307
rect 1479 301 1483 305
rect 1487 301 1489 305
rect 1479 299 1489 301
rect 1493 305 1503 307
rect 1493 301 1495 305
rect 1499 301 1503 305
rect 1493 299 1503 301
rect 1505 305 1515 307
rect 1505 301 1509 305
rect 1513 301 1515 305
rect 1505 299 1515 301
rect 1091 214 1101 216
rect 1091 210 1093 214
rect 1097 210 1101 214
rect 1091 208 1101 210
rect 1103 214 1113 216
rect 1103 210 1107 214
rect 1111 210 1113 214
rect 1103 208 1113 210
rect 1117 214 1127 216
rect 1117 210 1119 214
rect 1123 210 1127 214
rect 1117 208 1127 210
rect 1130 214 1142 216
rect 1130 210 1134 214
rect 1138 210 1142 214
rect 1130 208 1142 210
rect 1145 214 1155 216
rect 1145 210 1149 214
rect 1153 210 1155 214
rect 1145 208 1155 210
rect 1159 214 1169 216
rect 1159 210 1161 214
rect 1165 210 1169 214
rect 1159 208 1169 210
rect 1171 214 1181 216
rect 1171 210 1175 214
rect 1179 210 1181 214
rect 1171 208 1181 210
rect 1194 214 1204 216
rect 1194 210 1196 214
rect 1200 210 1204 214
rect 1194 208 1204 210
rect 1207 214 1219 216
rect 1207 210 1211 214
rect 1215 210 1219 214
rect 1207 208 1219 210
rect 1222 214 1234 216
rect 1222 210 1226 214
rect 1230 210 1234 214
rect 1222 208 1234 210
rect 1237 214 1249 216
rect 1237 210 1241 214
rect 1245 210 1249 214
rect 1237 208 1249 210
rect 1252 214 1262 216
rect 1252 210 1256 214
rect 1260 210 1262 214
rect 1252 208 1262 210
rect 1266 214 1276 216
rect 1266 210 1268 214
rect 1272 210 1276 214
rect 1266 208 1276 210
rect 1278 214 1288 216
rect 1278 210 1282 214
rect 1286 210 1288 214
rect 1278 208 1288 210
rect 759 206 769 208
rect 759 202 761 206
rect 765 202 769 206
rect 759 200 769 202
rect 771 206 781 208
rect 771 202 775 206
rect 779 202 781 206
rect 771 200 781 202
rect 785 206 795 208
rect 785 202 787 206
rect 791 202 795 206
rect 785 200 795 202
rect 798 206 810 208
rect 798 202 802 206
rect 806 202 810 206
rect 798 200 810 202
rect 813 206 823 208
rect 813 202 817 206
rect 821 202 823 206
rect 813 200 823 202
rect 827 206 837 208
rect 827 202 829 206
rect 833 202 837 206
rect 827 200 837 202
rect 839 206 849 208
rect 839 202 843 206
rect 847 202 849 206
rect 839 200 849 202
rect 866 206 876 208
rect 866 202 868 206
rect 872 202 876 206
rect 866 200 876 202
rect 879 206 891 208
rect 879 202 883 206
rect 887 202 891 206
rect 879 200 891 202
rect 894 206 906 208
rect 894 202 898 206
rect 902 202 906 206
rect 894 200 906 202
rect 909 206 919 208
rect 909 202 913 206
rect 917 202 919 206
rect 909 200 919 202
rect 923 206 933 208
rect 923 202 925 206
rect 929 202 933 206
rect 923 200 933 202
rect 935 206 945 208
rect 935 202 939 206
rect 943 202 945 206
rect 935 200 945 202
rect 414 193 424 195
rect 414 189 416 193
rect 420 189 424 193
rect 414 187 424 189
rect 426 193 436 195
rect 426 189 430 193
rect 434 189 436 193
rect 426 187 436 189
rect 440 193 450 195
rect 440 189 442 193
rect 446 189 450 193
rect 440 187 450 189
rect 453 193 465 195
rect 453 189 457 193
rect 461 189 465 193
rect 453 187 465 189
rect 468 193 478 195
rect 468 189 472 193
rect 476 189 478 193
rect 468 187 478 189
rect 482 193 492 195
rect 482 189 484 193
rect 488 189 492 193
rect 482 187 492 189
rect 494 193 504 195
rect 494 189 498 193
rect 502 189 504 193
rect 494 187 504 189
rect 517 193 527 195
rect 517 189 519 193
rect 523 189 527 193
rect 517 187 527 189
rect 530 193 542 195
rect 530 189 534 193
rect 538 189 542 193
rect 530 187 542 189
rect 545 193 555 195
rect 545 189 549 193
rect 553 189 555 193
rect 545 187 555 189
rect 559 193 569 195
rect 559 189 561 193
rect 565 189 569 193
rect 559 187 569 189
rect 571 193 581 195
rect 571 189 575 193
rect 579 189 581 193
rect 571 187 581 189
rect 68 150 78 152
rect 68 146 70 150
rect 74 146 78 150
rect 68 144 78 146
rect 80 150 90 152
rect 80 146 84 150
rect 88 146 90 150
rect 80 144 90 146
rect 94 150 104 152
rect 94 146 96 150
rect 100 146 104 150
rect 94 144 104 146
rect 107 150 119 152
rect 107 146 111 150
rect 115 146 119 150
rect 107 144 119 146
rect 122 150 132 152
rect 122 146 126 150
rect 130 146 132 150
rect 122 144 132 146
rect 136 150 146 152
rect 136 146 138 150
rect 142 146 146 150
rect 136 144 146 146
rect 148 150 158 152
rect 148 146 152 150
rect 156 146 158 150
rect 148 144 158 146
rect 1473 141 1483 143
rect 1473 137 1475 141
rect 1479 137 1483 141
rect 1473 135 1483 137
rect 1486 141 1498 143
rect 1486 137 1490 141
rect 1494 137 1498 141
rect 1486 135 1498 137
rect 1501 141 1513 143
rect 1501 137 1505 141
rect 1509 137 1513 141
rect 1501 135 1513 137
rect 1516 141 1528 143
rect 1516 137 1520 141
rect 1524 137 1528 141
rect 1516 135 1528 137
rect 1531 141 1541 143
rect 1531 137 1535 141
rect 1539 137 1541 141
rect 1531 135 1541 137
rect 1545 141 1555 143
rect 1545 137 1547 141
rect 1551 137 1555 141
rect 1545 135 1555 137
rect 1557 141 1567 143
rect 1557 137 1561 141
rect 1565 137 1567 141
rect 1557 135 1567 137
rect 1146 71 1156 73
rect 1146 67 1148 71
rect 1152 67 1156 71
rect 1146 65 1156 67
rect 1159 71 1171 73
rect 1159 67 1163 71
rect 1167 67 1171 71
rect 1159 65 1171 67
rect 1174 71 1184 73
rect 1174 67 1178 71
rect 1182 67 1184 71
rect 1174 65 1184 67
rect 802 63 812 65
rect 444 58 454 60
rect 98 55 108 57
rect 98 51 100 55
rect 104 51 108 55
rect 98 49 108 51
rect 111 55 123 57
rect 111 51 115 55
rect 119 51 123 55
rect 111 49 123 51
rect 126 55 136 57
rect 126 51 130 55
rect 134 51 136 55
rect 444 54 446 58
rect 450 54 454 58
rect 444 52 454 54
rect 457 58 469 60
rect 457 54 461 58
rect 465 54 469 58
rect 457 52 469 54
rect 472 58 482 60
rect 472 54 476 58
rect 480 54 482 58
rect 802 59 804 63
rect 808 59 812 63
rect 802 57 812 59
rect 815 63 827 65
rect 815 59 819 63
rect 823 59 827 63
rect 815 57 827 59
rect 830 63 840 65
rect 830 59 834 63
rect 838 59 840 63
rect 830 57 840 59
rect 472 52 482 54
rect 126 49 136 51
rect 31 16 41 18
rect 31 12 33 16
rect 37 12 41 16
rect 31 10 41 12
rect 44 16 56 18
rect 44 12 48 16
rect 52 12 56 16
rect 44 10 56 12
rect 59 16 69 18
rect 166 20 176 22
rect 59 12 63 16
rect 67 12 69 16
rect 59 10 69 12
rect 166 16 168 20
rect 172 16 176 20
rect 166 14 176 16
rect 179 20 191 22
rect 179 16 183 20
rect 187 16 191 20
rect 179 14 191 16
rect 194 20 204 22
rect 194 16 198 20
rect 202 16 204 20
rect 377 19 387 21
rect 194 14 204 16
rect 377 15 379 19
rect 383 15 387 19
rect 377 13 387 15
rect 390 19 402 21
rect 390 15 394 19
rect 398 15 402 19
rect 390 13 402 15
rect 405 19 415 21
rect 512 23 522 25
rect 405 15 409 19
rect 413 15 415 19
rect 405 13 415 15
rect 239 11 249 13
rect 239 7 241 11
rect 245 7 249 11
rect 239 5 249 7
rect 251 11 261 13
rect 251 7 255 11
rect 259 7 261 11
rect 251 5 261 7
rect 512 19 514 23
rect 518 19 522 23
rect 512 17 522 19
rect 525 23 537 25
rect 525 19 529 23
rect 533 19 537 23
rect 525 17 537 19
rect 540 23 550 25
rect 735 24 745 26
rect 540 19 544 23
rect 548 19 550 23
rect 735 20 737 24
rect 741 20 745 24
rect 540 17 550 19
rect 735 18 745 20
rect 748 24 760 26
rect 748 20 752 24
rect 756 20 760 24
rect 748 18 760 20
rect 763 24 773 26
rect 870 28 880 30
rect 763 20 767 24
rect 771 20 773 24
rect 763 18 773 20
rect 585 14 595 16
rect 585 10 587 14
rect 591 10 595 14
rect 585 8 595 10
rect 597 14 607 16
rect 597 10 601 14
rect 605 10 607 14
rect 597 8 607 10
rect 870 24 872 28
rect 876 24 880 28
rect 870 22 880 24
rect 883 28 895 30
rect 883 24 887 28
rect 891 24 895 28
rect 883 22 895 24
rect 898 28 908 30
rect 1079 32 1089 34
rect 898 24 902 28
rect 906 24 908 28
rect 1079 28 1081 32
rect 1085 28 1089 32
rect 1079 26 1089 28
rect 1092 32 1104 34
rect 1092 28 1096 32
rect 1100 28 1104 32
rect 1092 26 1104 28
rect 1107 32 1117 34
rect 1214 36 1224 38
rect 1107 28 1111 32
rect 1115 28 1117 32
rect 1107 26 1117 28
rect 898 22 908 24
rect 943 19 953 21
rect 943 15 945 19
rect 949 15 953 19
rect 943 13 953 15
rect 955 19 965 21
rect 955 15 959 19
rect 963 15 965 19
rect 955 13 965 15
rect 1214 32 1216 36
rect 1220 32 1224 36
rect 1214 30 1224 32
rect 1227 36 1239 38
rect 1227 32 1231 36
rect 1235 32 1239 36
rect 1227 30 1239 32
rect 1242 36 1252 38
rect 1242 32 1246 36
rect 1250 32 1252 36
rect 1242 30 1252 32
rect 1287 27 1297 29
rect 1287 23 1289 27
rect 1293 23 1297 27
rect 1287 21 1297 23
rect 1299 27 1309 29
rect 1299 23 1303 27
rect 1307 23 1309 27
rect 1299 21 1309 23
rect 98 -28 108 -26
rect 98 -32 100 -28
rect 104 -32 108 -28
rect 98 -34 108 -32
rect 111 -28 123 -26
rect 111 -32 115 -28
rect 119 -32 123 -28
rect 111 -34 123 -32
rect 126 -28 136 -26
rect 444 -25 454 -23
rect 126 -32 130 -28
rect 134 -32 136 -28
rect 444 -29 446 -25
rect 450 -29 454 -25
rect 444 -31 454 -29
rect 457 -25 469 -23
rect 457 -29 461 -25
rect 465 -29 469 -25
rect 457 -31 469 -29
rect 472 -25 482 -23
rect 1146 -12 1156 -10
rect 802 -20 812 -18
rect 802 -24 804 -20
rect 808 -24 812 -20
rect 472 -29 476 -25
rect 480 -29 482 -25
rect 802 -26 812 -24
rect 815 -20 827 -18
rect 815 -24 819 -20
rect 823 -24 827 -20
rect 815 -26 827 -24
rect 830 -20 840 -18
rect 1146 -16 1148 -12
rect 1152 -16 1156 -12
rect 1146 -18 1156 -16
rect 1159 -12 1171 -10
rect 1159 -16 1163 -12
rect 1167 -16 1171 -12
rect 1159 -18 1171 -16
rect 1174 -12 1184 -10
rect 1174 -16 1178 -12
rect 1182 -16 1184 -12
rect 1174 -18 1184 -16
rect 830 -24 834 -20
rect 838 -24 840 -20
rect 830 -26 840 -24
rect 472 -31 482 -29
rect 126 -34 136 -32
rect 76 -130 86 -128
rect 76 -134 78 -130
rect 82 -134 86 -130
rect 76 -136 86 -134
rect 88 -130 98 -128
rect 88 -134 92 -130
rect 96 -134 98 -130
rect 88 -136 98 -134
rect 102 -130 112 -128
rect 102 -134 104 -130
rect 108 -134 112 -130
rect 102 -136 112 -134
rect 115 -130 127 -128
rect 115 -134 119 -130
rect 123 -134 127 -130
rect 115 -136 127 -134
rect 130 -130 140 -128
rect 130 -134 134 -130
rect 138 -134 140 -130
rect 130 -136 140 -134
rect 144 -130 154 -128
rect 144 -134 146 -130
rect 150 -134 154 -130
rect 144 -136 154 -134
rect 156 -130 166 -128
rect 156 -134 160 -130
rect 164 -134 166 -130
rect 156 -136 166 -134
rect 1077 -157 1087 -155
rect 731 -159 741 -157
rect 731 -163 733 -159
rect 737 -163 741 -159
rect 731 -165 741 -163
rect 743 -159 753 -157
rect 743 -163 747 -159
rect 751 -163 753 -159
rect 743 -165 753 -163
rect 757 -159 767 -157
rect 757 -163 759 -159
rect 763 -163 767 -159
rect 757 -165 767 -163
rect 770 -159 782 -157
rect 770 -163 774 -159
rect 778 -163 782 -159
rect 770 -165 782 -163
rect 785 -159 795 -157
rect 785 -163 789 -159
rect 793 -163 795 -159
rect 785 -165 795 -163
rect 799 -159 809 -157
rect 799 -163 801 -159
rect 805 -163 809 -159
rect 799 -165 809 -163
rect 811 -159 821 -157
rect 811 -163 815 -159
rect 819 -163 821 -159
rect 811 -165 821 -163
rect 838 -159 848 -157
rect 838 -163 840 -159
rect 844 -163 848 -159
rect 838 -165 848 -163
rect 851 -159 863 -157
rect 851 -163 855 -159
rect 859 -163 863 -159
rect 851 -165 863 -163
rect 866 -159 878 -157
rect 866 -163 870 -159
rect 874 -163 878 -159
rect 866 -165 878 -163
rect 881 -159 891 -157
rect 881 -163 885 -159
rect 889 -163 891 -159
rect 881 -165 891 -163
rect 895 -159 905 -157
rect 895 -163 897 -159
rect 901 -163 905 -159
rect 895 -165 905 -163
rect 907 -159 917 -157
rect 907 -163 911 -159
rect 915 -163 917 -159
rect 1077 -161 1079 -157
rect 1083 -161 1087 -157
rect 1077 -163 1087 -161
rect 1089 -157 1099 -155
rect 1089 -161 1093 -157
rect 1097 -161 1099 -157
rect 1089 -163 1099 -161
rect 1103 -157 1113 -155
rect 1103 -161 1105 -157
rect 1109 -161 1113 -157
rect 1103 -163 1113 -161
rect 1116 -157 1128 -155
rect 1116 -161 1120 -157
rect 1124 -161 1128 -157
rect 1116 -163 1128 -161
rect 1131 -157 1141 -155
rect 1131 -161 1135 -157
rect 1139 -161 1141 -157
rect 1131 -163 1141 -161
rect 1145 -157 1155 -155
rect 1145 -161 1147 -157
rect 1151 -161 1155 -157
rect 1145 -163 1155 -161
rect 1157 -157 1167 -155
rect 1157 -161 1161 -157
rect 1165 -161 1167 -157
rect 1157 -163 1167 -161
rect 1180 -157 1190 -155
rect 1180 -161 1182 -157
rect 1186 -161 1190 -157
rect 1180 -163 1190 -161
rect 1193 -157 1205 -155
rect 1193 -161 1197 -157
rect 1201 -161 1205 -157
rect 1193 -163 1205 -161
rect 1208 -157 1220 -155
rect 1208 -161 1212 -157
rect 1216 -161 1220 -157
rect 1208 -163 1220 -161
rect 1223 -157 1235 -155
rect 1223 -161 1227 -157
rect 1231 -161 1235 -157
rect 1223 -163 1235 -161
rect 1238 -157 1248 -155
rect 1238 -161 1242 -157
rect 1246 -161 1248 -157
rect 1238 -163 1248 -161
rect 1252 -157 1262 -155
rect 1252 -161 1254 -157
rect 1258 -161 1262 -157
rect 1252 -163 1262 -161
rect 1264 -157 1274 -155
rect 1264 -161 1268 -157
rect 1272 -161 1274 -157
rect 1264 -163 1274 -161
rect 907 -165 917 -163
rect 406 -174 416 -172
rect 406 -178 408 -174
rect 412 -178 416 -174
rect 406 -180 416 -178
rect 418 -174 428 -172
rect 418 -178 422 -174
rect 426 -178 428 -174
rect 418 -180 428 -178
rect 432 -174 442 -172
rect 432 -178 434 -174
rect 438 -178 442 -174
rect 432 -180 442 -178
rect 445 -174 457 -172
rect 445 -178 449 -174
rect 453 -178 457 -174
rect 445 -180 457 -178
rect 460 -174 470 -172
rect 460 -178 464 -174
rect 468 -178 470 -174
rect 460 -180 470 -178
rect 474 -174 484 -172
rect 474 -178 476 -174
rect 480 -178 484 -174
rect 474 -180 484 -178
rect 486 -174 496 -172
rect 486 -178 490 -174
rect 494 -178 496 -174
rect 486 -180 496 -178
rect 509 -174 519 -172
rect 509 -178 511 -174
rect 515 -178 519 -174
rect 509 -180 519 -178
rect 522 -174 534 -172
rect 522 -178 526 -174
rect 530 -178 534 -174
rect 522 -180 534 -178
rect 537 -174 547 -172
rect 537 -178 541 -174
rect 545 -178 547 -174
rect 537 -180 547 -178
rect 551 -174 561 -172
rect 551 -178 553 -174
rect 557 -178 561 -174
rect 551 -180 561 -178
rect 563 -174 573 -172
rect 563 -178 567 -174
rect 571 -178 573 -174
rect 563 -180 573 -178
rect 1339 -358 1349 -356
rect 1339 -362 1341 -358
rect 1345 -362 1349 -358
rect 1339 -364 1349 -362
rect 1352 -364 1373 -356
rect 1376 -364 1399 -356
rect 1402 -364 1423 -356
rect 1426 -358 1436 -356
rect 1426 -362 1430 -358
rect 1434 -362 1436 -358
rect 1426 -364 1436 -362
rect 1440 -358 1450 -356
rect 1440 -362 1442 -358
rect 1446 -362 1450 -358
rect 1440 -364 1450 -362
rect 1452 -358 1462 -356
rect 1452 -362 1456 -358
rect 1460 -362 1462 -358
rect 1452 -364 1462 -362
<< metal1 >>
rect -30 137 -26 370
rect -30 133 -28 137
rect -30 -5 -26 133
rect -13 120 -9 372
rect 316 294 320 370
rect 333 294 337 370
rect 674 294 678 370
rect 691 294 695 369
rect 1018 294 1022 370
rect 1035 294 1039 369
rect 1439 319 1443 406
rect 1392 315 1399 319
rect 1403 315 1423 319
rect 1427 315 1449 319
rect 1453 315 1477 319
rect 1481 315 1495 319
rect 1499 315 1509 319
rect 1513 315 1517 319
rect 1394 305 1398 315
rect 1495 305 1499 315
rect 173 290 175 294
rect 1341 290 1472 294
rect 66 160 70 164
rect 74 160 84 164
rect 88 160 101 164
rect 105 160 120 164
rect 124 160 138 164
rect 142 160 152 164
rect 156 160 158 164
rect 70 150 74 160
rect 96 150 100 160
rect 126 150 130 160
rect 138 150 142 160
rect 68 133 73 137
rect 84 121 88 146
rect 111 137 115 146
rect 98 133 103 137
rect 111 133 130 137
rect 99 129 103 133
rect 126 129 130 133
rect 152 131 156 146
rect 173 131 177 290
rect 316 180 320 290
rect 316 176 318 180
rect 99 125 114 129
rect 126 125 142 129
rect 152 127 177 131
rect 286 130 288 134
rect -13 116 -11 120
rect 68 116 74 120
rect 84 117 99 121
rect -30 -9 -28 -5
rect -30 -160 -26 -9
rect -13 -13 -9 116
rect 84 110 88 117
rect 126 110 130 125
rect 152 110 156 127
rect 70 98 74 106
rect 96 98 100 106
rect 138 98 142 106
rect 68 94 70 98
rect 74 94 85 98
rect 89 94 101 98
rect 105 94 122 98
rect 126 94 138 98
rect 142 94 153 98
rect 157 94 158 98
rect 98 65 105 69
rect 109 65 124 69
rect 128 65 136 69
rect 100 55 104 65
rect 130 55 134 65
rect 115 42 119 51
rect 115 38 134 42
rect 21 34 96 38
rect 130 34 134 38
rect 21 -5 26 34
rect 92 30 118 34
rect 130 30 150 34
rect 166 30 173 34
rect 177 30 192 34
rect 196 30 237 34
rect 29 26 38 30
rect 42 26 57 30
rect 61 26 66 30
rect 33 16 37 26
rect 63 16 67 26
rect 83 22 103 26
rect 48 3 52 12
rect 48 -1 67 3
rect 63 -5 67 -1
rect 83 -5 87 22
rect 130 15 134 30
rect 100 3 104 11
rect 98 -1 105 3
rect 109 -1 126 3
rect 130 -1 134 3
rect 146 -1 150 30
rect 168 20 172 30
rect 198 20 202 30
rect 233 25 237 30
rect 233 21 241 25
rect 245 21 255 25
rect 259 21 263 25
rect 183 7 187 16
rect 241 11 245 21
rect 183 3 202 7
rect 198 -1 202 3
rect 255 0 259 7
rect 286 0 290 130
rect 146 -5 186 -1
rect 198 -5 245 -1
rect 255 -4 290 0
rect 12 -9 51 -5
rect 63 -9 87 -5
rect -13 -17 -11 -13
rect 12 -17 36 -13
rect -13 -143 -9 -17
rect 23 -44 28 -17
rect 63 -24 67 -9
rect 33 -36 37 -28
rect 31 -40 38 -36
rect 42 -40 59 -36
rect 63 -40 68 -36
rect 23 -48 78 -44
rect 73 -57 78 -48
rect 83 -49 87 -9
rect 146 -13 171 -9
rect 99 -18 105 -14
rect 109 -18 124 -14
rect 128 -18 136 -14
rect 100 -28 104 -18
rect 130 -28 134 -18
rect 115 -41 119 -32
rect 115 -45 134 -41
rect 130 -49 134 -45
rect 146 -49 150 -13
rect 198 -20 202 -5
rect 255 -11 259 -4
rect 241 -23 245 -15
rect 168 -32 172 -24
rect 235 -27 241 -23
rect 245 -27 256 -23
rect 260 -27 263 -23
rect 168 -36 173 -32
rect 177 -36 194 -32
rect 198 -40 202 -32
rect 235 -40 239 -27
rect 198 -44 239 -40
rect 83 -53 118 -49
rect 130 -53 150 -49
rect 73 -61 103 -57
rect 130 -68 134 -53
rect 100 -80 104 -72
rect 100 -84 105 -80
rect 109 -84 126 -80
rect 130 -84 134 -80
rect 115 -88 119 -84
rect 74 -120 78 -116
rect 82 -120 92 -116
rect 96 -120 109 -116
rect 113 -120 128 -116
rect 132 -120 146 -116
rect 150 -120 160 -116
rect 164 -120 166 -116
rect 78 -130 82 -120
rect 104 -130 108 -120
rect 134 -130 138 -120
rect 146 -130 150 -120
rect -13 -147 -11 -143
rect 76 -147 81 -143
rect -30 -164 -28 -160
rect -30 -190 -26 -164
rect -13 -188 -9 -147
rect 92 -159 96 -134
rect 119 -143 123 -134
rect 106 -147 111 -143
rect 119 -147 138 -143
rect 107 -151 111 -147
rect 134 -151 138 -147
rect 160 -149 164 -134
rect 107 -155 122 -151
rect 134 -155 150 -151
rect 160 -153 184 -149
rect 76 -164 82 -160
rect 92 -163 107 -159
rect 92 -170 96 -163
rect 134 -170 138 -155
rect 160 -170 164 -153
rect 78 -182 82 -174
rect 104 -182 108 -174
rect 146 -182 150 -174
rect 76 -186 78 -182
rect 82 -186 93 -182
rect 97 -186 109 -182
rect 113 -186 130 -182
rect 134 -186 146 -182
rect 150 -186 161 -182
rect 165 -186 166 -182
rect 180 -390 184 -153
rect 286 -275 290 -4
rect 316 -2 320 176
rect 333 163 337 290
rect 674 287 678 290
rect 691 287 695 290
rect 1018 287 1022 290
rect 1035 287 1039 290
rect 591 283 593 287
rect 1339 283 1448 287
rect 1483 284 1487 301
rect 1509 286 1513 301
rect 413 203 416 207
rect 420 203 430 207
rect 434 203 447 207
rect 451 203 466 207
rect 470 203 484 207
rect 488 203 498 207
rect 502 203 524 207
rect 528 203 543 207
rect 547 203 561 207
rect 565 203 575 207
rect 579 203 581 207
rect 416 193 420 203
rect 442 193 446 203
rect 472 193 476 203
rect 484 193 488 203
rect 519 193 523 203
rect 549 193 553 203
rect 561 193 565 203
rect 414 176 419 180
rect 430 164 434 189
rect 457 180 461 189
rect 444 176 449 180
rect 457 176 476 180
rect 445 172 449 176
rect 472 172 476 176
rect 498 172 502 189
rect 534 180 538 189
rect 534 176 553 180
rect 549 172 553 176
rect 575 174 579 189
rect 591 174 595 283
rect 445 168 460 172
rect 472 168 488 172
rect 498 168 537 172
rect 549 168 565 172
rect 575 170 595 174
rect 674 193 678 283
rect 674 189 676 193
rect 333 159 335 163
rect 414 159 420 163
rect 430 160 445 164
rect 316 -6 318 -2
rect 316 -204 320 -6
rect 333 -10 337 159
rect 430 153 434 160
rect 472 153 476 168
rect 498 153 502 168
rect 549 153 553 168
rect 575 153 579 170
rect 416 141 420 149
rect 442 141 446 149
rect 484 141 488 149
rect 519 141 523 149
rect 561 141 565 149
rect 414 137 416 141
rect 420 137 431 141
rect 435 137 447 141
rect 451 137 468 141
rect 472 137 484 141
rect 488 137 499 141
rect 503 137 524 141
rect 528 137 545 141
rect 549 137 561 141
rect 565 137 576 141
rect 580 137 585 141
rect 632 120 635 124
rect 444 68 451 72
rect 455 68 470 72
rect 474 68 482 72
rect 446 58 450 68
rect 476 58 480 68
rect 461 45 465 54
rect 461 41 480 45
rect 367 37 442 41
rect 476 37 480 41
rect 367 -2 372 37
rect 438 33 464 37
rect 476 33 496 37
rect 512 33 519 37
rect 523 33 538 37
rect 542 33 583 37
rect 375 29 384 33
rect 388 29 403 33
rect 407 29 412 33
rect 379 19 383 29
rect 409 19 413 29
rect 429 25 449 29
rect 394 6 398 15
rect 394 2 413 6
rect 409 -2 413 2
rect 429 -2 433 25
rect 476 18 480 33
rect 446 6 450 14
rect 444 2 451 6
rect 455 2 472 6
rect 476 2 480 6
rect 492 2 496 33
rect 514 23 518 33
rect 544 23 548 33
rect 579 28 583 33
rect 579 24 587 28
rect 591 24 601 28
rect 605 24 609 28
rect 529 10 533 19
rect 587 14 591 24
rect 529 6 548 10
rect 544 2 548 6
rect 601 3 605 10
rect 632 3 637 120
rect 492 -2 532 2
rect 544 -2 591 2
rect 601 -1 637 3
rect 358 -6 397 -2
rect 409 -6 433 -2
rect 333 -14 335 -10
rect 358 -14 382 -10
rect 333 -187 337 -14
rect 369 -41 374 -14
rect 409 -21 413 -6
rect 379 -33 383 -25
rect 377 -37 384 -33
rect 388 -37 405 -33
rect 409 -37 414 -33
rect 369 -45 424 -41
rect 419 -54 424 -45
rect 429 -46 433 -6
rect 492 -10 517 -6
rect 445 -15 451 -11
rect 455 -15 470 -11
rect 474 -15 482 -11
rect 446 -25 450 -15
rect 476 -25 480 -15
rect 461 -38 465 -29
rect 461 -42 480 -38
rect 476 -46 480 -42
rect 492 -46 496 -10
rect 544 -17 548 -2
rect 601 -8 605 -1
rect 587 -20 591 -12
rect 514 -29 518 -21
rect 581 -24 587 -20
rect 591 -24 602 -20
rect 606 -24 609 -20
rect 514 -33 519 -29
rect 523 -33 540 -29
rect 544 -37 548 -29
rect 581 -37 585 -24
rect 544 -41 585 -37
rect 429 -50 464 -46
rect 476 -50 496 -46
rect 419 -58 449 -54
rect 476 -65 480 -50
rect 446 -77 450 -69
rect 446 -81 451 -77
rect 455 -81 472 -77
rect 476 -81 480 -77
rect 461 -85 465 -81
rect 405 -164 408 -160
rect 412 -164 422 -160
rect 426 -164 439 -160
rect 443 -164 458 -160
rect 462 -164 476 -160
rect 480 -164 490 -160
rect 494 -164 516 -160
rect 520 -164 535 -160
rect 539 -164 553 -160
rect 557 -164 567 -160
rect 571 -164 572 -160
rect 408 -174 412 -164
rect 434 -174 438 -164
rect 464 -174 468 -164
rect 476 -174 480 -164
rect 511 -174 515 -164
rect 541 -174 545 -164
rect 553 -174 557 -164
rect 333 -191 335 -187
rect 406 -191 411 -187
rect 316 -208 318 -204
rect 316 -230 320 -208
rect 333 -230 337 -191
rect 422 -203 426 -178
rect 449 -187 453 -178
rect 436 -191 441 -187
rect 449 -191 468 -187
rect 437 -195 441 -191
rect 464 -195 468 -191
rect 490 -195 494 -178
rect 526 -187 530 -178
rect 526 -191 545 -187
rect 541 -195 545 -191
rect 567 -193 571 -178
rect 437 -199 452 -195
rect 464 -199 480 -195
rect 490 -199 529 -195
rect 541 -199 557 -195
rect 567 -197 594 -193
rect 406 -208 412 -204
rect 422 -207 437 -203
rect 422 -214 426 -207
rect 464 -214 468 -199
rect 490 -214 494 -199
rect 541 -214 545 -199
rect 567 -214 571 -197
rect 408 -226 412 -218
rect 434 -226 438 -218
rect 476 -226 480 -218
rect 511 -226 515 -218
rect 553 -226 557 -218
rect 406 -230 408 -226
rect 412 -230 423 -226
rect 427 -230 439 -226
rect 443 -230 460 -226
rect 464 -230 476 -226
rect 480 -230 491 -226
rect 495 -230 516 -226
rect 520 -230 537 -226
rect 541 -230 553 -226
rect 557 -230 568 -226
rect 572 -230 575 -226
rect 286 -279 292 -275
rect 590 -383 594 -197
rect 632 -266 637 -1
rect 674 3 678 189
rect 691 176 695 283
rect 1018 280 1022 283
rect 1035 280 1039 283
rect 1458 280 1499 284
rect 1509 282 1517 286
rect 960 276 962 280
rect 1337 276 1422 280
rect 758 216 761 220
rect 765 216 775 220
rect 779 216 792 220
rect 796 216 811 220
rect 815 216 829 220
rect 833 216 843 220
rect 847 216 873 220
rect 877 216 907 220
rect 911 216 925 220
rect 929 216 939 220
rect 943 216 945 220
rect 761 206 765 216
rect 787 206 791 216
rect 817 206 821 216
rect 829 206 833 216
rect 868 206 872 216
rect 913 206 917 216
rect 759 189 764 193
rect 775 177 779 202
rect 802 193 806 202
rect 789 189 794 193
rect 802 189 821 193
rect 790 185 794 189
rect 817 185 821 189
rect 843 187 847 202
rect 883 195 887 202
rect 925 206 929 216
rect 898 195 902 202
rect 853 191 872 195
rect 883 191 917 195
rect 853 187 857 191
rect 790 181 805 185
rect 817 181 833 185
rect 843 183 857 187
rect 913 184 917 191
rect 939 186 943 202
rect 960 186 964 276
rect 691 172 693 176
rect 759 172 765 176
rect 775 173 790 177
rect 674 -1 676 3
rect 674 -189 678 -1
rect 691 -5 695 172
rect 775 166 779 173
rect 817 166 821 181
rect 843 166 847 183
rect 913 180 929 184
rect 939 182 964 186
rect 1018 201 1022 276
rect 1018 197 1020 201
rect 862 170 902 174
rect 913 165 917 180
rect 939 165 943 182
rect 761 154 765 162
rect 787 154 791 162
rect 829 154 833 162
rect 759 150 761 154
rect 765 150 776 154
rect 780 150 792 154
rect 796 150 813 154
rect 817 150 829 154
rect 833 150 844 154
rect 848 153 862 154
rect 868 153 872 161
rect 925 153 929 161
rect 848 150 873 153
rect 857 149 873 150
rect 877 149 909 153
rect 913 149 925 153
rect 929 149 940 153
rect 944 149 945 153
rect 902 126 906 142
rect 979 111 981 115
rect 802 73 809 77
rect 813 73 828 77
rect 832 73 840 77
rect 804 63 808 73
rect 834 63 838 73
rect 819 50 823 59
rect 819 46 838 50
rect 725 42 800 46
rect 834 42 838 46
rect 725 3 730 42
rect 796 38 822 42
rect 834 38 854 42
rect 870 38 877 42
rect 881 38 896 42
rect 900 38 941 42
rect 733 34 742 38
rect 746 34 761 38
rect 765 34 770 38
rect 737 24 741 34
rect 767 24 771 34
rect 787 30 807 34
rect 752 11 756 20
rect 752 7 771 11
rect 767 3 771 7
rect 787 3 791 30
rect 834 23 838 38
rect 804 11 808 19
rect 802 7 809 11
rect 813 7 830 11
rect 834 7 838 11
rect 850 7 854 38
rect 872 28 876 38
rect 902 28 906 38
rect 937 33 941 38
rect 937 29 945 33
rect 949 29 959 33
rect 963 29 967 33
rect 887 15 891 24
rect 945 19 949 29
rect 887 11 906 15
rect 902 7 906 11
rect 959 8 963 15
rect 979 8 983 111
rect 850 3 890 7
rect 902 3 949 7
rect 959 4 983 8
rect 716 -1 755 3
rect 767 -1 791 3
rect 691 -9 693 -5
rect 716 -9 740 -5
rect 691 -172 695 -9
rect 727 -36 732 -9
rect 767 -16 771 -1
rect 737 -28 741 -20
rect 735 -32 742 -28
rect 746 -32 763 -28
rect 767 -32 772 -28
rect 727 -40 782 -36
rect 777 -49 782 -40
rect 787 -41 791 -1
rect 850 -5 875 -1
rect 803 -10 809 -6
rect 813 -10 828 -6
rect 832 -10 840 -6
rect 804 -20 808 -10
rect 834 -20 838 -10
rect 819 -33 823 -24
rect 819 -37 838 -33
rect 834 -41 838 -37
rect 850 -41 854 -5
rect 902 -12 906 3
rect 959 -3 963 4
rect 945 -15 949 -7
rect 872 -24 876 -16
rect 939 -19 945 -15
rect 949 -19 960 -15
rect 964 -19 967 -15
rect 872 -28 877 -24
rect 881 -28 898 -24
rect 902 -32 906 -24
rect 939 -32 943 -19
rect 902 -36 943 -32
rect 787 -45 822 -41
rect 834 -45 854 -41
rect 777 -53 807 -49
rect 834 -60 838 -45
rect 804 -72 808 -64
rect 804 -76 809 -72
rect 813 -76 830 -72
rect 834 -76 838 -72
rect 819 -80 823 -76
rect 730 -149 733 -145
rect 737 -149 747 -145
rect 751 -149 764 -145
rect 768 -149 783 -145
rect 787 -149 801 -145
rect 805 -149 815 -145
rect 819 -149 845 -145
rect 849 -149 879 -145
rect 883 -149 897 -145
rect 901 -149 911 -145
rect 915 -149 919 -145
rect 733 -159 737 -149
rect 759 -159 763 -149
rect 789 -159 793 -149
rect 801 -159 805 -149
rect 840 -159 844 -149
rect 885 -159 889 -149
rect 691 -176 693 -172
rect 731 -176 736 -172
rect 674 -193 676 -189
rect 674 -245 678 -193
rect 691 -236 695 -176
rect 747 -188 751 -163
rect 774 -172 778 -163
rect 761 -176 766 -172
rect 774 -176 793 -172
rect 762 -180 766 -176
rect 789 -180 793 -176
rect 815 -178 819 -163
rect 855 -170 859 -163
rect 897 -159 901 -149
rect 870 -170 874 -163
rect 825 -174 844 -170
rect 855 -174 889 -170
rect 825 -178 829 -174
rect 762 -184 777 -180
rect 789 -184 805 -180
rect 815 -182 829 -178
rect 885 -181 889 -174
rect 911 -179 915 -163
rect 731 -193 737 -189
rect 747 -192 762 -188
rect 747 -199 751 -192
rect 789 -199 793 -184
rect 815 -199 819 -182
rect 885 -185 901 -181
rect 911 -183 948 -179
rect 834 -195 874 -191
rect 885 -200 889 -185
rect 911 -200 915 -183
rect 733 -211 737 -203
rect 759 -211 763 -203
rect 801 -211 805 -203
rect 731 -215 733 -211
rect 737 -215 748 -211
rect 752 -215 764 -211
rect 768 -215 785 -211
rect 789 -215 801 -211
rect 805 -215 816 -211
rect 820 -212 834 -211
rect 840 -212 844 -204
rect 897 -212 901 -204
rect 820 -215 845 -212
rect 829 -216 845 -215
rect 849 -216 881 -212
rect 885 -216 897 -212
rect 901 -216 912 -212
rect 916 -216 918 -212
rect 632 -270 635 -266
rect 878 -273 882 -257
rect 944 -376 948 -183
rect 979 -256 983 4
rect 1018 11 1022 197
rect 1035 184 1039 276
rect 1458 273 1462 280
rect 1326 269 1398 273
rect 1408 269 1462 273
rect 1091 224 1093 228
rect 1097 224 1107 228
rect 1111 224 1124 228
rect 1128 224 1143 228
rect 1147 224 1161 228
rect 1165 224 1175 228
rect 1179 224 1201 228
rect 1205 224 1250 228
rect 1254 224 1268 228
rect 1272 224 1282 228
rect 1286 224 1288 228
rect 1093 214 1097 224
rect 1119 214 1123 224
rect 1149 214 1153 224
rect 1161 214 1165 224
rect 1196 214 1200 224
rect 1256 214 1260 224
rect 1091 197 1096 201
rect 1107 185 1111 210
rect 1134 201 1138 210
rect 1121 197 1126 201
rect 1134 197 1153 201
rect 1122 193 1126 197
rect 1149 193 1153 197
rect 1175 195 1179 210
rect 1211 203 1215 210
rect 1226 203 1230 210
rect 1268 214 1272 224
rect 1241 203 1245 210
rect 1183 199 1200 203
rect 1211 199 1260 203
rect 1183 195 1187 199
rect 1122 189 1137 193
rect 1149 189 1165 193
rect 1175 191 1187 195
rect 1256 192 1260 199
rect 1282 194 1286 210
rect 1326 194 1330 269
rect 1408 264 1412 269
rect 1432 264 1436 269
rect 1458 264 1462 269
rect 1483 264 1487 280
rect 1509 264 1513 282
rect 1394 252 1398 260
rect 1418 252 1422 260
rect 1444 252 1448 260
rect 1468 252 1472 260
rect 1495 252 1499 260
rect 1392 248 1399 252
rect 1403 248 1423 252
rect 1427 248 1449 252
rect 1453 248 1479 252
rect 1483 248 1495 252
rect 1499 248 1510 252
rect 1514 248 1515 252
rect 1035 180 1037 184
rect 1091 180 1097 184
rect 1107 181 1122 185
rect 1018 7 1020 11
rect 1018 -187 1022 7
rect 1035 3 1039 180
rect 1107 174 1111 181
rect 1149 174 1153 189
rect 1175 174 1179 191
rect 1256 188 1272 192
rect 1282 190 1330 194
rect 1256 173 1260 188
rect 1282 173 1286 190
rect 1093 162 1097 170
rect 1119 162 1123 170
rect 1161 162 1165 170
rect 1091 158 1093 162
rect 1097 158 1108 162
rect 1112 158 1124 162
rect 1128 158 1145 162
rect 1149 158 1161 162
rect 1165 158 1176 162
rect 1180 161 1192 162
rect 1196 161 1200 169
rect 1268 161 1272 169
rect 1411 166 1512 170
rect 1180 158 1201 161
rect 1189 157 1201 158
rect 1205 157 1252 161
rect 1256 157 1268 161
rect 1272 157 1283 161
rect 1287 157 1288 161
rect 1234 126 1238 140
rect 1244 117 1248 140
rect 1146 81 1153 85
rect 1157 81 1172 85
rect 1176 81 1318 85
rect 1148 71 1152 81
rect 1178 71 1182 81
rect 1163 58 1167 67
rect 1314 62 1318 81
rect 1411 62 1415 166
rect 1508 155 1512 166
rect 1473 151 1480 155
rect 1484 151 1529 155
rect 1533 151 1547 155
rect 1551 151 1561 155
rect 1565 151 1569 155
rect 1475 141 1479 151
rect 1535 141 1539 151
rect 1490 130 1494 137
rect 1505 130 1509 137
rect 1547 141 1551 151
rect 1520 130 1524 137
rect 1471 126 1479 130
rect 1490 126 1539 130
rect 1471 119 1494 123
rect 1535 119 1539 126
rect 1561 121 1565 137
rect 1471 112 1509 116
rect 1535 115 1551 119
rect 1561 117 1569 121
rect 1471 105 1524 109
rect 1535 100 1539 115
rect 1561 100 1565 117
rect 1475 88 1479 96
rect 1547 88 1551 96
rect 1473 84 1480 88
rect 1484 84 1531 88
rect 1535 84 1547 88
rect 1551 84 1562 88
rect 1566 84 1567 88
rect 1314 58 1415 62
rect 1163 54 1182 58
rect 1069 50 1144 54
rect 1178 50 1182 54
rect 1069 11 1074 50
rect 1140 46 1166 50
rect 1178 46 1198 50
rect 1214 46 1221 50
rect 1225 46 1240 50
rect 1244 46 1285 50
rect 1077 42 1086 46
rect 1090 42 1105 46
rect 1109 42 1114 46
rect 1081 32 1085 42
rect 1111 32 1115 42
rect 1131 38 1151 42
rect 1096 19 1100 28
rect 1096 15 1115 19
rect 1111 11 1115 15
rect 1131 11 1135 38
rect 1178 31 1182 46
rect 1148 19 1152 27
rect 1146 15 1153 19
rect 1157 15 1174 19
rect 1178 15 1182 19
rect 1194 15 1198 46
rect 1216 36 1220 46
rect 1246 36 1250 46
rect 1281 41 1285 46
rect 1281 37 1289 41
rect 1293 37 1303 41
rect 1307 37 1311 41
rect 1231 23 1235 32
rect 1289 27 1293 37
rect 1231 19 1250 23
rect 1246 15 1250 19
rect 1303 16 1307 23
rect 1194 11 1234 15
rect 1246 11 1293 15
rect 1303 12 1313 16
rect 1060 7 1099 11
rect 1111 7 1135 11
rect 1035 -1 1037 3
rect 1060 -1 1084 3
rect 1035 -170 1039 -1
rect 1071 -28 1076 -1
rect 1111 -8 1115 7
rect 1081 -20 1085 -12
rect 1079 -24 1086 -20
rect 1090 -24 1107 -20
rect 1111 -24 1116 -20
rect 1071 -32 1126 -28
rect 1121 -41 1126 -32
rect 1131 -33 1135 7
rect 1194 3 1219 7
rect 1147 -2 1153 2
rect 1157 -2 1172 2
rect 1176 -2 1184 2
rect 1148 -12 1152 -2
rect 1178 -12 1182 -2
rect 1163 -25 1167 -16
rect 1163 -29 1182 -25
rect 1178 -33 1182 -29
rect 1194 -33 1198 3
rect 1246 -4 1250 11
rect 1303 5 1307 12
rect 1289 -7 1293 1
rect 1216 -16 1220 -8
rect 1283 -11 1289 -7
rect 1293 -11 1304 -7
rect 1308 -11 1311 -7
rect 1216 -20 1221 -16
rect 1225 -20 1242 -16
rect 1246 -24 1250 -16
rect 1283 -24 1287 -11
rect 1246 -28 1287 -24
rect 1131 -37 1166 -33
rect 1178 -37 1198 -33
rect 1121 -45 1151 -41
rect 1178 -52 1182 -37
rect 1148 -64 1152 -56
rect 1148 -68 1153 -64
rect 1157 -68 1174 -64
rect 1178 -68 1182 -64
rect 1163 -72 1167 -68
rect 1411 -143 1415 58
rect 1075 -147 1079 -143
rect 1083 -147 1093 -143
rect 1097 -147 1110 -143
rect 1114 -147 1129 -143
rect 1133 -147 1147 -143
rect 1151 -147 1161 -143
rect 1165 -147 1187 -143
rect 1191 -147 1236 -143
rect 1240 -147 1254 -143
rect 1258 -147 1268 -143
rect 1272 -147 1415 -143
rect 1079 -157 1083 -147
rect 1105 -157 1109 -147
rect 1135 -157 1139 -147
rect 1147 -157 1151 -147
rect 1182 -157 1186 -147
rect 1242 -157 1246 -147
rect 1035 -174 1037 -170
rect 1077 -174 1082 -170
rect 1018 -191 1020 -187
rect 1018 -213 1022 -191
rect 1035 -213 1039 -174
rect 1093 -186 1097 -161
rect 1120 -170 1124 -161
rect 1107 -174 1112 -170
rect 1120 -174 1139 -170
rect 1108 -178 1112 -174
rect 1135 -178 1139 -174
rect 1161 -176 1165 -161
rect 1197 -168 1201 -161
rect 1212 -168 1216 -161
rect 1254 -157 1258 -147
rect 1227 -168 1231 -161
rect 1169 -172 1186 -168
rect 1197 -172 1246 -168
rect 1169 -176 1173 -172
rect 1108 -182 1123 -178
rect 1135 -182 1151 -178
rect 1161 -180 1173 -176
rect 1242 -179 1246 -172
rect 1268 -177 1272 -161
rect 1077 -191 1083 -187
rect 1093 -190 1108 -186
rect 1093 -197 1097 -190
rect 1135 -197 1139 -182
rect 1161 -197 1165 -180
rect 1242 -183 1258 -179
rect 1268 -181 1302 -177
rect 1242 -198 1246 -183
rect 1268 -198 1272 -181
rect 1079 -209 1083 -201
rect 1105 -209 1109 -201
rect 1147 -209 1151 -201
rect 1077 -213 1079 -209
rect 1083 -213 1094 -209
rect 1098 -213 1110 -209
rect 1114 -213 1131 -209
rect 1135 -213 1147 -209
rect 1151 -213 1162 -209
rect 1166 -210 1178 -209
rect 1182 -210 1186 -202
rect 1254 -210 1258 -202
rect 1166 -213 1187 -210
rect 1175 -214 1187 -213
rect 1191 -214 1238 -210
rect 1242 -214 1254 -210
rect 1258 -214 1269 -210
rect 1273 -214 1274 -210
rect 979 -260 981 -256
rect 1220 -264 1224 -247
rect 1235 -273 1239 -247
rect 1297 -369 1302 -181
rect 1411 -344 1415 -147
rect 1337 -348 1346 -344
rect 1350 -348 1370 -344
rect 1374 -348 1396 -344
rect 1400 -348 1424 -344
rect 1428 -348 1442 -344
rect 1446 -348 1456 -344
rect 1460 -348 1464 -344
rect 1341 -358 1345 -348
rect 1442 -358 1446 -348
rect 1297 -373 1419 -369
rect 944 -380 1395 -376
rect 1430 -379 1434 -362
rect 1456 -377 1460 -362
rect 1405 -383 1446 -379
rect 1456 -381 1464 -377
rect 590 -387 1369 -383
rect 1405 -390 1409 -383
rect 180 -394 1345 -390
rect 1355 -394 1409 -390
rect 1355 -399 1359 -394
rect 1379 -399 1383 -394
rect 1405 -399 1409 -394
rect 1430 -399 1434 -383
rect 1456 -399 1460 -381
rect 1341 -411 1345 -403
rect 1365 -411 1369 -403
rect 1391 -411 1395 -403
rect 1415 -411 1419 -403
rect 1442 -411 1446 -403
rect 1339 -415 1346 -411
rect 1350 -415 1370 -411
rect 1374 -415 1396 -411
rect 1400 -415 1426 -411
rect 1430 -415 1442 -411
rect 1446 -415 1457 -411
rect 1461 -415 1464 -411
rect 1385 -451 1389 -415
<< metal2 >>
rect 1373 315 1388 319
rect 1373 228 1377 315
rect 1519 248 1600 252
rect 1073 224 1087 228
rect 1292 224 1377 228
rect 1073 220 1077 224
rect 720 216 754 220
rect 949 216 1077 220
rect 720 207 724 216
rect 277 203 409 207
rect 585 203 724 207
rect 277 164 281 203
rect 1100 197 1117 201
rect 768 189 785 193
rect 423 176 440 180
rect 162 160 281 164
rect 1071 158 1087 162
rect 740 150 755 154
rect 1071 153 1075 158
rect 1292 157 1357 161
rect 740 141 744 150
rect 949 149 1075 153
rect 269 137 410 141
rect 589 137 744 141
rect 77 133 94 137
rect 269 98 273 137
rect 162 94 273 98
rect 1353 88 1357 157
rect 1373 155 1377 224
rect 1373 151 1469 155
rect 1596 88 1600 248
rect 1116 81 1142 85
rect 1353 84 1469 88
rect 1571 84 1600 88
rect 1116 77 1120 81
rect 772 73 798 77
rect 844 73 1120 77
rect 772 72 776 73
rect 414 69 440 72
rect 68 65 94 69
rect 140 68 440 69
rect 486 68 776 72
rect 140 65 418 68
rect 68 30 72 65
rect 139 38 214 42
rect 70 26 80 30
rect 76 -14 80 26
rect 139 3 143 38
rect 138 -1 143 3
rect 155 30 162 34
rect 155 -14 159 30
rect 76 -18 95 -14
rect 140 -18 159 -14
rect 210 -32 214 38
rect 414 33 418 65
rect 485 41 560 45
rect 416 29 426 33
rect 422 -11 426 29
rect 485 6 489 41
rect 484 2 489 6
rect 501 33 508 37
rect 501 -11 505 33
rect 422 -15 441 -11
rect 486 -15 505 -11
rect 556 -29 560 41
rect 772 38 776 68
rect 843 46 918 50
rect 1116 46 1120 73
rect 1187 54 1262 58
rect 774 34 784 38
rect 780 -6 784 34
rect 843 11 847 46
rect 842 7 847 11
rect 859 38 866 42
rect 859 -6 863 38
rect 780 -10 799 -6
rect 844 -10 863 -6
rect 914 -24 918 46
rect 1118 42 1128 46
rect 1124 2 1128 42
rect 1187 19 1191 54
rect 1186 15 1191 19
rect 1203 46 1210 50
rect 1203 2 1207 46
rect 1124 -2 1143 2
rect 1188 -2 1207 2
rect 1258 -16 1262 54
rect 1210 -20 1212 -16
rect 1254 -20 1262 -16
rect 1120 -24 1130 -20
rect 866 -28 868 -24
rect 910 -28 918 -24
rect 162 -36 164 -32
rect 206 -36 214 -32
rect 508 -33 510 -29
rect 552 -33 560 -29
rect 776 -32 786 -28
rect 72 -40 82 -36
rect 78 -80 82 -40
rect 162 -80 166 -36
rect 418 -37 428 -33
rect 424 -77 428 -37
rect 508 -76 512 -33
rect 782 -71 786 -32
rect 754 -72 786 -71
rect 866 -70 870 -28
rect 1126 -61 1130 -24
rect 1106 -64 1130 -61
rect 1210 -61 1214 -20
rect 1376 -61 1380 84
rect 1210 -64 1380 -61
rect 1106 -65 1144 -64
rect 1106 -70 1110 -65
rect 1126 -68 1144 -65
rect 1186 -65 1380 -64
rect 1186 -68 1214 -65
rect 866 -72 1110 -70
rect 754 -75 800 -72
rect 754 -76 758 -75
rect 782 -76 800 -75
rect 842 -74 1110 -72
rect 842 -76 870 -74
rect 508 -77 758 -76
rect 401 -80 442 -77
rect 78 -84 96 -80
rect 138 -81 442 -80
rect 484 -80 758 -77
rect 484 -81 512 -80
rect 138 -84 405 -81
rect 170 -120 394 -116
rect 85 -147 102 -143
rect 390 -160 394 -120
rect 1055 -145 1070 -143
rect 705 -149 726 -145
rect 923 -147 1070 -145
rect 923 -149 1059 -147
rect 705 -160 709 -149
rect 390 -164 401 -160
rect 576 -164 709 -160
rect 740 -176 757 -172
rect 1086 -174 1103 -170
rect 170 -186 302 -182
rect 298 -226 302 -186
rect 415 -191 432 -187
rect 710 -215 727 -211
rect 1057 -212 1073 -209
rect 710 -226 714 -215
rect 922 -213 1073 -212
rect 1376 -210 1380 -65
rect 922 -216 1061 -213
rect 1278 -214 1380 -210
rect 298 -230 402 -226
rect 579 -230 714 -226
rect 1278 -411 1282 -214
rect 1278 -415 1335 -411
<< ntransistor >>
rect 1402 258 1405 266
rect 1426 258 1429 266
rect 1452 258 1455 266
rect 1476 258 1479 266
rect 1503 258 1505 266
rect 424 147 426 155
rect 450 147 453 155
rect 465 147 468 155
rect 492 147 494 155
rect 769 160 771 168
rect 795 160 798 168
rect 810 160 813 168
rect 837 160 839 168
rect 1101 168 1103 176
rect 1127 168 1130 176
rect 1142 168 1145 176
rect 1169 168 1171 176
rect 876 159 879 167
rect 891 159 894 167
rect 906 159 909 167
rect 933 159 935 167
rect 1204 167 1207 175
rect 1219 167 1222 175
rect 1234 167 1237 175
rect 1249 167 1252 175
rect 1276 167 1278 175
rect 527 147 530 155
rect 542 147 545 155
rect 569 147 571 155
rect 78 104 80 112
rect 104 104 107 112
rect 119 104 122 112
rect 146 104 148 112
rect 108 9 111 17
rect 123 9 126 17
rect 249 -17 251 -9
rect 454 12 457 20
rect 469 12 472 20
rect 41 -30 44 -22
rect 56 -30 59 -22
rect 176 -26 179 -18
rect 191 -26 194 -18
rect 812 17 815 25
rect 827 17 830 25
rect 595 -14 597 -6
rect 1156 25 1159 33
rect 1171 25 1174 33
rect 953 -9 955 -1
rect 1483 94 1486 102
rect 1498 94 1501 102
rect 1513 94 1516 102
rect 1528 94 1531 102
rect 1555 94 1557 102
rect 1297 -1 1299 7
rect 387 -27 390 -19
rect 402 -27 405 -19
rect 522 -23 525 -15
rect 537 -23 540 -15
rect 745 -22 748 -14
rect 760 -22 763 -14
rect 880 -18 883 -10
rect 895 -18 898 -10
rect 1089 -14 1092 -6
rect 1104 -14 1107 -6
rect 1224 -10 1227 -2
rect 1239 -10 1242 -2
rect 1156 -58 1159 -50
rect 1171 -58 1174 -50
rect 108 -74 111 -66
rect 123 -74 126 -66
rect 454 -71 457 -63
rect 469 -71 472 -63
rect 812 -66 815 -58
rect 827 -66 830 -58
rect 86 -176 88 -168
rect 112 -176 115 -168
rect 127 -176 130 -168
rect 154 -176 156 -168
rect 416 -220 418 -212
rect 442 -220 445 -212
rect 457 -220 460 -212
rect 484 -220 486 -212
rect 741 -205 743 -197
rect 767 -205 770 -197
rect 782 -205 785 -197
rect 809 -205 811 -197
rect 848 -206 851 -198
rect 863 -206 866 -198
rect 878 -206 881 -198
rect 905 -206 907 -198
rect 1087 -203 1089 -195
rect 1113 -203 1116 -195
rect 1128 -203 1131 -195
rect 1155 -203 1157 -195
rect 1190 -204 1193 -196
rect 1205 -204 1208 -196
rect 1220 -204 1223 -196
rect 1235 -204 1238 -196
rect 1262 -204 1264 -196
rect 519 -220 522 -212
rect 534 -220 537 -212
rect 561 -220 563 -212
rect 1349 -405 1352 -397
rect 1373 -405 1376 -397
rect 1399 -405 1402 -397
rect 1423 -405 1426 -397
rect 1450 -405 1452 -397
<< ptransistor >>
rect 1402 299 1405 307
rect 1426 299 1429 307
rect 1452 299 1455 307
rect 1476 299 1479 307
rect 1503 299 1505 307
rect 1101 208 1103 216
rect 1127 208 1130 216
rect 1142 208 1145 216
rect 1169 208 1171 216
rect 1204 208 1207 216
rect 1219 208 1222 216
rect 1234 208 1237 216
rect 1249 208 1252 216
rect 1276 208 1278 216
rect 769 200 771 208
rect 795 200 798 208
rect 810 200 813 208
rect 837 200 839 208
rect 876 200 879 208
rect 891 200 894 208
rect 906 200 909 208
rect 933 200 935 208
rect 424 187 426 195
rect 450 187 453 195
rect 465 187 468 195
rect 492 187 494 195
rect 527 187 530 195
rect 542 187 545 195
rect 569 187 571 195
rect 78 144 80 152
rect 104 144 107 152
rect 119 144 122 152
rect 146 144 148 152
rect 1483 135 1486 143
rect 1498 135 1501 143
rect 1513 135 1516 143
rect 1528 135 1531 143
rect 1555 135 1557 143
rect 1156 65 1159 73
rect 1171 65 1174 73
rect 108 49 111 57
rect 123 49 126 57
rect 454 52 457 60
rect 469 52 472 60
rect 812 57 815 65
rect 827 57 830 65
rect 41 10 44 18
rect 56 10 59 18
rect 176 14 179 22
rect 191 14 194 22
rect 387 13 390 21
rect 402 13 405 21
rect 249 5 251 13
rect 522 17 525 25
rect 537 17 540 25
rect 745 18 748 26
rect 760 18 763 26
rect 595 8 597 16
rect 880 22 883 30
rect 895 22 898 30
rect 1089 26 1092 34
rect 1104 26 1107 34
rect 953 13 955 21
rect 1224 30 1227 38
rect 1239 30 1242 38
rect 1297 21 1299 29
rect 108 -34 111 -26
rect 123 -34 126 -26
rect 454 -31 457 -23
rect 469 -31 472 -23
rect 812 -26 815 -18
rect 827 -26 830 -18
rect 1156 -18 1159 -10
rect 1171 -18 1174 -10
rect 86 -136 88 -128
rect 112 -136 115 -128
rect 127 -136 130 -128
rect 154 -136 156 -128
rect 741 -165 743 -157
rect 767 -165 770 -157
rect 782 -165 785 -157
rect 809 -165 811 -157
rect 848 -165 851 -157
rect 863 -165 866 -157
rect 878 -165 881 -157
rect 905 -165 907 -157
rect 1087 -163 1089 -155
rect 1113 -163 1116 -155
rect 1128 -163 1131 -155
rect 1155 -163 1157 -155
rect 1190 -163 1193 -155
rect 1205 -163 1208 -155
rect 1220 -163 1223 -155
rect 1235 -163 1238 -155
rect 1262 -163 1264 -155
rect 416 -180 418 -172
rect 442 -180 445 -172
rect 457 -180 460 -172
rect 484 -180 486 -172
rect 519 -180 522 -172
rect 534 -180 537 -172
rect 561 -180 563 -172
rect 1349 -364 1352 -356
rect 1373 -364 1376 -356
rect 1399 -364 1402 -356
rect 1423 -364 1426 -356
rect 1450 -364 1452 -356
<< polycontact >>
rect 175 290 179 294
rect 1337 290 1341 294
rect 593 283 597 287
rect 1335 283 1339 287
rect 962 276 966 280
rect 1333 276 1337 280
rect 1398 269 1402 273
rect 1422 276 1426 280
rect 1448 283 1452 287
rect 1472 290 1476 294
rect 1499 280 1503 284
rect 676 189 680 193
rect 755 189 759 193
rect 318 176 322 180
rect 410 176 414 180
rect 335 159 339 163
rect 410 159 414 163
rect 420 159 424 163
rect 460 168 464 172
rect 488 168 492 172
rect 445 160 449 164
rect 537 168 541 172
rect 565 168 569 172
rect -28 133 -24 137
rect 64 133 68 137
rect -11 116 -7 120
rect 64 116 68 120
rect 74 116 78 120
rect 114 125 118 129
rect 142 125 146 129
rect 99 117 103 121
rect 693 172 697 176
rect 755 172 759 176
rect 765 172 769 176
rect 805 181 809 185
rect 833 181 837 185
rect 790 173 794 177
rect 872 191 876 195
rect 902 170 906 174
rect 929 180 933 184
rect 1020 197 1024 201
rect 1087 197 1091 201
rect 1037 180 1041 184
rect 1087 180 1091 184
rect 1097 180 1101 184
rect 1137 189 1141 193
rect 1165 189 1169 193
rect 1122 181 1126 185
rect 1200 199 1204 203
rect 1272 188 1276 192
rect 902 142 906 146
rect 1234 140 1238 144
rect 1244 140 1248 144
rect 288 130 292 134
rect 1467 126 1471 130
rect 1479 126 1483 130
rect 635 120 639 124
rect 902 122 906 126
rect 1234 122 1238 126
rect 1467 119 1471 123
rect 981 111 985 115
rect 1244 113 1248 117
rect 1467 112 1471 116
rect 1467 105 1471 109
rect 1494 119 1498 123
rect 1509 112 1513 116
rect 1524 105 1528 109
rect 1551 115 1555 119
rect 118 30 122 34
rect 103 22 107 26
rect 464 33 468 37
rect 1166 46 1170 50
rect 822 38 826 42
rect 1151 38 1155 42
rect 449 25 453 29
rect -28 -9 -24 -5
rect 8 -9 12 -5
rect 51 -9 55 -5
rect 807 30 811 34
rect 186 -5 190 -1
rect 245 -5 249 -1
rect -11 -17 -7 -13
rect 8 -17 12 -13
rect 36 -17 40 -13
rect 171 -13 175 -9
rect 318 -6 322 -2
rect 354 -6 358 -2
rect 397 -6 401 -2
rect 532 -2 536 2
rect 591 -2 595 2
rect 335 -14 339 -10
rect 354 -14 358 -10
rect 382 -14 386 -10
rect 517 -10 521 -6
rect 676 -1 680 3
rect 712 -1 716 3
rect 755 -1 759 3
rect 890 3 894 7
rect 949 3 953 7
rect 693 -9 697 -5
rect 712 -9 716 -5
rect 740 -9 744 -5
rect 875 -5 879 -1
rect 1020 7 1024 11
rect 1056 7 1060 11
rect 1099 7 1103 11
rect 1234 11 1238 15
rect 1293 11 1297 15
rect 1037 -1 1041 3
rect 1056 -1 1060 3
rect 1084 -1 1088 3
rect 1219 3 1223 7
rect 1313 12 1317 16
rect 118 -53 122 -49
rect 103 -61 107 -57
rect 464 -50 468 -46
rect 1166 -37 1170 -33
rect 822 -45 826 -41
rect 1151 -45 1155 -41
rect 449 -58 453 -54
rect 807 -53 811 -49
rect -11 -147 -7 -143
rect 72 -147 76 -143
rect -28 -164 -24 -160
rect 72 -164 76 -160
rect 82 -164 86 -160
rect 122 -155 126 -151
rect 150 -155 154 -151
rect 107 -163 111 -159
rect 693 -176 697 -172
rect 727 -176 731 -172
rect 335 -191 339 -187
rect 402 -191 406 -187
rect 318 -208 322 -204
rect 402 -208 406 -204
rect 412 -208 416 -204
rect 452 -199 456 -195
rect 480 -199 484 -195
rect 437 -207 441 -203
rect 529 -199 533 -195
rect 557 -199 561 -195
rect 676 -193 680 -189
rect 727 -193 731 -189
rect 737 -193 741 -189
rect 777 -184 781 -180
rect 805 -184 809 -180
rect 762 -192 766 -188
rect 844 -174 848 -170
rect 874 -195 878 -191
rect 901 -185 905 -181
rect 1037 -174 1041 -170
rect 1073 -174 1077 -170
rect 1020 -191 1024 -187
rect 1073 -191 1077 -187
rect 1083 -191 1087 -187
rect 1123 -182 1127 -178
rect 1151 -182 1155 -178
rect 1108 -190 1112 -186
rect 1186 -172 1190 -168
rect 1258 -183 1262 -179
rect 878 -257 882 -253
rect 1220 -247 1224 -243
rect 1235 -247 1239 -243
rect 981 -260 985 -256
rect 635 -270 639 -266
rect 1220 -268 1224 -264
rect 292 -279 296 -275
rect 878 -277 882 -273
rect 1235 -277 1239 -273
rect 1345 -394 1349 -390
rect 1369 -387 1373 -383
rect 1395 -380 1399 -376
rect 1419 -373 1423 -369
rect 1446 -383 1450 -379
<< ndcontact >>
rect 1394 260 1398 264
rect 1408 260 1412 264
rect 1418 260 1422 264
rect 1432 260 1436 264
rect 1444 260 1448 264
rect 1458 260 1462 264
rect 1468 260 1472 264
rect 1483 260 1487 264
rect 1495 260 1499 264
rect 1509 260 1513 264
rect 416 149 420 153
rect 430 149 434 153
rect 442 149 446 153
rect 472 149 476 153
rect 484 149 488 153
rect 498 149 502 153
rect 761 162 765 166
rect 775 162 779 166
rect 787 162 791 166
rect 817 162 821 166
rect 829 162 833 166
rect 1093 170 1097 174
rect 1107 170 1111 174
rect 1119 170 1123 174
rect 1149 170 1153 174
rect 1161 170 1165 174
rect 1175 170 1179 174
rect 1196 169 1200 173
rect 843 162 847 166
rect 868 161 872 165
rect 913 161 917 165
rect 925 161 929 165
rect 1256 169 1260 173
rect 1268 169 1272 173
rect 1282 169 1286 173
rect 939 161 943 165
rect 519 149 523 153
rect 549 149 553 153
rect 561 149 565 153
rect 575 149 579 153
rect 70 106 74 110
rect 84 106 88 110
rect 96 106 100 110
rect 126 106 130 110
rect 138 106 142 110
rect 152 106 156 110
rect 100 11 104 15
rect 130 11 134 15
rect 446 14 450 18
rect 241 -15 245 -11
rect 476 14 480 18
rect 804 19 808 23
rect 255 -15 259 -11
rect 33 -28 37 -24
rect 63 -28 67 -24
rect 168 -24 172 -20
rect 834 19 838 23
rect 1148 27 1152 31
rect 587 -12 591 -8
rect 601 -12 605 -8
rect 1178 27 1182 31
rect 945 -7 949 -3
rect 959 -7 963 -3
rect 1475 96 1479 100
rect 1535 96 1539 100
rect 1547 96 1551 100
rect 1561 96 1565 100
rect 1289 1 1293 5
rect 1303 1 1307 5
rect 198 -24 202 -20
rect 379 -25 383 -21
rect 409 -25 413 -21
rect 514 -21 518 -17
rect 544 -21 548 -17
rect 737 -20 741 -16
rect 767 -20 771 -16
rect 872 -16 876 -12
rect 902 -16 906 -12
rect 1081 -12 1085 -8
rect 1111 -12 1115 -8
rect 1216 -8 1220 -4
rect 1246 -8 1250 -4
rect 1148 -56 1152 -52
rect 1178 -56 1182 -52
rect 100 -72 104 -68
rect 130 -72 134 -68
rect 446 -69 450 -65
rect 476 -69 480 -65
rect 804 -64 808 -60
rect 834 -64 838 -60
rect 78 -174 82 -170
rect 92 -174 96 -170
rect 104 -174 108 -170
rect 134 -174 138 -170
rect 146 -174 150 -170
rect 160 -174 164 -170
rect 408 -218 412 -214
rect 422 -218 426 -214
rect 434 -218 438 -214
rect 464 -218 468 -214
rect 476 -218 480 -214
rect 490 -218 494 -214
rect 733 -203 737 -199
rect 747 -203 751 -199
rect 759 -203 763 -199
rect 789 -203 793 -199
rect 801 -203 805 -199
rect 815 -203 819 -199
rect 840 -204 844 -200
rect 885 -204 889 -200
rect 897 -204 901 -200
rect 911 -204 915 -200
rect 1079 -201 1083 -197
rect 1093 -201 1097 -197
rect 1105 -201 1109 -197
rect 1135 -201 1139 -197
rect 1147 -201 1151 -197
rect 1161 -201 1165 -197
rect 1182 -202 1186 -198
rect 1242 -202 1246 -198
rect 1254 -202 1258 -198
rect 1268 -202 1272 -198
rect 511 -218 515 -214
rect 541 -218 545 -214
rect 553 -218 557 -214
rect 567 -218 571 -214
rect 1341 -403 1345 -399
rect 1355 -403 1359 -399
rect 1365 -403 1369 -399
rect 1379 -403 1383 -399
rect 1391 -403 1395 -399
rect 1405 -403 1409 -399
rect 1415 -403 1419 -399
rect 1430 -403 1434 -399
rect 1442 -403 1446 -399
rect 1456 -403 1460 -399
<< pdcontact >>
rect 1394 301 1398 305
rect 1483 301 1487 305
rect 1495 301 1499 305
rect 1509 301 1513 305
rect 1093 210 1097 214
rect 1107 210 1111 214
rect 1119 210 1123 214
rect 1134 210 1138 214
rect 1149 210 1153 214
rect 1161 210 1165 214
rect 1175 210 1179 214
rect 1196 210 1200 214
rect 1211 210 1215 214
rect 1226 210 1230 214
rect 1241 210 1245 214
rect 1256 210 1260 214
rect 1268 210 1272 214
rect 1282 210 1286 214
rect 761 202 765 206
rect 775 202 779 206
rect 787 202 791 206
rect 802 202 806 206
rect 817 202 821 206
rect 829 202 833 206
rect 843 202 847 206
rect 868 202 872 206
rect 883 202 887 206
rect 898 202 902 206
rect 913 202 917 206
rect 925 202 929 206
rect 939 202 943 206
rect 416 189 420 193
rect 430 189 434 193
rect 442 189 446 193
rect 457 189 461 193
rect 472 189 476 193
rect 484 189 488 193
rect 498 189 502 193
rect 519 189 523 193
rect 534 189 538 193
rect 549 189 553 193
rect 561 189 565 193
rect 575 189 579 193
rect 70 146 74 150
rect 84 146 88 150
rect 96 146 100 150
rect 111 146 115 150
rect 126 146 130 150
rect 138 146 142 150
rect 152 146 156 150
rect 1475 137 1479 141
rect 1490 137 1494 141
rect 1505 137 1509 141
rect 1520 137 1524 141
rect 1535 137 1539 141
rect 1547 137 1551 141
rect 1561 137 1565 141
rect 1148 67 1152 71
rect 1163 67 1167 71
rect 1178 67 1182 71
rect 100 51 104 55
rect 115 51 119 55
rect 130 51 134 55
rect 446 54 450 58
rect 461 54 465 58
rect 476 54 480 58
rect 804 59 808 63
rect 819 59 823 63
rect 834 59 838 63
rect 33 12 37 16
rect 48 12 52 16
rect 63 12 67 16
rect 168 16 172 20
rect 183 16 187 20
rect 198 16 202 20
rect 379 15 383 19
rect 394 15 398 19
rect 409 15 413 19
rect 241 7 245 11
rect 255 7 259 11
rect 514 19 518 23
rect 529 19 533 23
rect 544 19 548 23
rect 737 20 741 24
rect 752 20 756 24
rect 767 20 771 24
rect 587 10 591 14
rect 601 10 605 14
rect 872 24 876 28
rect 887 24 891 28
rect 902 24 906 28
rect 1081 28 1085 32
rect 1096 28 1100 32
rect 1111 28 1115 32
rect 945 15 949 19
rect 959 15 963 19
rect 1216 32 1220 36
rect 1231 32 1235 36
rect 1246 32 1250 36
rect 1289 23 1293 27
rect 1303 23 1307 27
rect 100 -32 104 -28
rect 115 -32 119 -28
rect 130 -32 134 -28
rect 446 -29 450 -25
rect 461 -29 465 -25
rect 804 -24 808 -20
rect 476 -29 480 -25
rect 819 -24 823 -20
rect 1148 -16 1152 -12
rect 1163 -16 1167 -12
rect 1178 -16 1182 -12
rect 834 -24 838 -20
rect 78 -134 82 -130
rect 92 -134 96 -130
rect 104 -134 108 -130
rect 119 -134 123 -130
rect 134 -134 138 -130
rect 146 -134 150 -130
rect 160 -134 164 -130
rect 733 -163 737 -159
rect 747 -163 751 -159
rect 759 -163 763 -159
rect 774 -163 778 -159
rect 789 -163 793 -159
rect 801 -163 805 -159
rect 815 -163 819 -159
rect 840 -163 844 -159
rect 855 -163 859 -159
rect 870 -163 874 -159
rect 885 -163 889 -159
rect 897 -163 901 -159
rect 911 -163 915 -159
rect 1079 -161 1083 -157
rect 1093 -161 1097 -157
rect 1105 -161 1109 -157
rect 1120 -161 1124 -157
rect 1135 -161 1139 -157
rect 1147 -161 1151 -157
rect 1161 -161 1165 -157
rect 1182 -161 1186 -157
rect 1197 -161 1201 -157
rect 1212 -161 1216 -157
rect 1227 -161 1231 -157
rect 1242 -161 1246 -157
rect 1254 -161 1258 -157
rect 1268 -161 1272 -157
rect 408 -178 412 -174
rect 422 -178 426 -174
rect 434 -178 438 -174
rect 449 -178 453 -174
rect 464 -178 468 -174
rect 476 -178 480 -174
rect 490 -178 494 -174
rect 511 -178 515 -174
rect 526 -178 530 -174
rect 541 -178 545 -174
rect 553 -178 557 -174
rect 567 -178 571 -174
rect 1341 -362 1345 -358
rect 1430 -362 1434 -358
rect 1442 -362 1446 -358
rect 1456 -362 1460 -358
<< nbccdiffcontact >>
rect 1495 315 1499 319
rect 1093 224 1097 228
rect 1161 224 1165 228
rect 1268 224 1272 228
rect 761 216 765 220
rect 829 216 833 220
rect 925 216 929 220
rect 416 203 420 207
rect 484 203 488 207
rect 561 203 565 207
rect 70 160 74 164
rect 138 160 142 164
rect 1547 151 1551 155
rect 241 21 245 25
rect 587 24 591 28
rect 945 29 949 33
rect 1289 37 1293 41
rect 78 -120 82 -116
rect 146 -120 150 -116
rect 733 -149 737 -145
rect 801 -149 805 -145
rect 897 -149 901 -145
rect 1079 -147 1083 -143
rect 1147 -147 1151 -143
rect 1254 -147 1258 -143
rect 408 -164 412 -160
rect 476 -164 480 -160
rect 553 -164 557 -160
rect 1442 -348 1446 -344
<< m2contact >>
rect 1388 315 1392 319
rect 158 160 162 164
rect 73 133 77 137
rect 94 133 98 137
rect 158 94 162 98
rect 94 65 98 69
rect 136 65 140 69
rect 162 30 166 34
rect 66 26 70 30
rect 134 -1 138 3
rect 68 -40 72 -36
rect 95 -18 99 -14
rect 136 -18 140 -14
rect 164 -36 168 -32
rect 202 -36 206 -32
rect 96 -84 100 -80
rect 134 -84 138 -80
rect 166 -120 170 -116
rect 81 -147 85 -143
rect 102 -147 106 -143
rect 166 -186 170 -182
rect 409 203 413 207
rect 581 203 585 207
rect 419 176 423 180
rect 440 176 444 180
rect 410 137 414 141
rect 585 137 589 141
rect 440 68 444 72
rect 482 68 486 72
rect 508 33 512 37
rect 412 29 416 33
rect 480 2 484 6
rect 414 -37 418 -33
rect 441 -15 445 -11
rect 482 -15 486 -11
rect 510 -33 514 -29
rect 548 -33 552 -29
rect 442 -81 446 -77
rect 480 -81 484 -77
rect 401 -164 405 -160
rect 572 -164 576 -160
rect 411 -191 415 -187
rect 432 -191 436 -187
rect 402 -230 406 -226
rect 575 -230 579 -226
rect 754 216 758 220
rect 945 216 949 220
rect 764 189 768 193
rect 785 189 789 193
rect 755 150 759 154
rect 945 149 949 153
rect 798 73 802 77
rect 840 73 844 77
rect 866 38 870 42
rect 770 34 774 38
rect 838 7 842 11
rect 772 -32 776 -28
rect 799 -10 803 -6
rect 840 -10 844 -6
rect 868 -28 872 -24
rect 906 -28 910 -24
rect 800 -76 804 -72
rect 838 -76 842 -72
rect 726 -149 730 -145
rect 919 -149 923 -145
rect 736 -176 740 -172
rect 757 -176 761 -172
rect 727 -215 731 -211
rect 918 -216 922 -212
rect 1087 224 1091 228
rect 1288 224 1292 228
rect 1096 197 1100 201
rect 1117 197 1121 201
rect 1515 248 1519 252
rect 1087 158 1091 162
rect 1288 157 1292 161
rect 1142 81 1146 85
rect 1469 151 1473 155
rect 1469 84 1473 88
rect 1567 84 1571 88
rect 1210 46 1214 50
rect 1114 42 1118 46
rect 1182 15 1186 19
rect 1116 -24 1120 -20
rect 1143 -2 1147 2
rect 1184 -2 1188 2
rect 1212 -20 1216 -16
rect 1250 -20 1254 -16
rect 1144 -68 1148 -64
rect 1182 -68 1186 -64
rect 1070 -147 1075 -143
rect 1082 -174 1086 -170
rect 1103 -174 1107 -170
rect 1073 -213 1077 -209
rect 1274 -214 1278 -210
rect 1335 -415 1339 -411
<< psubstratepcontact >>
rect 1399 248 1403 252
rect 1423 248 1427 252
rect 1449 248 1453 252
rect 1479 248 1483 252
rect 1495 248 1499 252
rect 1510 248 1514 252
rect 416 137 420 141
rect 431 137 435 141
rect 447 137 451 141
rect 468 137 472 141
rect 484 137 488 141
rect 499 137 503 141
rect 761 150 765 154
rect 776 150 780 154
rect 792 150 796 154
rect 813 150 817 154
rect 829 150 833 154
rect 844 150 848 154
rect 873 149 877 153
rect 524 137 528 141
rect 545 137 549 141
rect 561 137 565 141
rect 576 137 580 141
rect 1093 158 1097 162
rect 1108 158 1112 162
rect 1124 158 1128 162
rect 1145 158 1149 162
rect 1161 158 1165 162
rect 1176 158 1180 162
rect 1201 157 1205 161
rect 909 149 913 153
rect 925 149 929 153
rect 940 149 944 153
rect 1252 157 1256 161
rect 1268 157 1272 161
rect 1283 157 1287 161
rect 70 94 74 98
rect 85 94 89 98
rect 101 94 105 98
rect 122 94 126 98
rect 138 94 142 98
rect 153 94 157 98
rect 105 -1 109 3
rect 126 -1 130 3
rect 451 2 455 6
rect 472 2 476 6
rect 809 7 813 11
rect 830 7 834 11
rect 1153 15 1157 19
rect 1174 15 1178 19
rect 1480 84 1484 88
rect 1531 84 1535 88
rect 1547 84 1551 88
rect 1562 84 1566 88
rect 241 -27 245 -23
rect 256 -27 260 -23
rect 587 -24 591 -20
rect 602 -24 606 -20
rect 945 -19 949 -15
rect 960 -19 964 -15
rect 1289 -11 1293 -7
rect 1304 -11 1308 -7
rect 1086 -24 1090 -20
rect 1107 -24 1111 -20
rect 38 -40 42 -36
rect 59 -40 63 -36
rect 173 -36 177 -32
rect 194 -36 198 -32
rect 384 -37 388 -33
rect 405 -37 409 -33
rect 519 -33 523 -29
rect 540 -33 544 -29
rect 742 -32 746 -28
rect 763 -32 767 -28
rect 877 -28 881 -24
rect 898 -28 902 -24
rect 1221 -20 1225 -16
rect 1242 -20 1246 -16
rect 1153 -68 1157 -64
rect 1174 -68 1178 -64
rect 809 -76 813 -72
rect 830 -76 834 -72
rect 105 -84 109 -80
rect 126 -84 130 -80
rect 451 -81 455 -77
rect 472 -81 476 -77
rect 78 -186 82 -182
rect 93 -186 97 -182
rect 109 -186 113 -182
rect 130 -186 134 -182
rect 146 -186 150 -182
rect 161 -186 165 -182
rect 408 -230 412 -226
rect 423 -230 427 -226
rect 439 -230 443 -226
rect 460 -230 464 -226
rect 476 -230 480 -226
rect 491 -230 495 -226
rect 733 -215 737 -211
rect 748 -215 752 -211
rect 764 -215 768 -211
rect 785 -215 789 -211
rect 801 -215 805 -211
rect 816 -215 820 -211
rect 845 -216 849 -212
rect 516 -230 520 -226
rect 537 -230 541 -226
rect 553 -230 557 -226
rect 568 -230 572 -226
rect 881 -216 885 -212
rect 897 -216 901 -212
rect 912 -216 916 -212
rect 1079 -213 1083 -209
rect 1094 -213 1098 -209
rect 1110 -213 1114 -209
rect 1131 -213 1135 -209
rect 1147 -213 1151 -209
rect 1162 -213 1166 -209
rect 1187 -214 1191 -210
rect 1238 -214 1242 -210
rect 1254 -214 1258 -210
rect 1269 -214 1273 -210
rect 1346 -415 1350 -411
rect 1370 -415 1374 -411
rect 1396 -415 1400 -411
rect 1426 -415 1430 -411
rect 1442 -415 1446 -411
rect 1457 -415 1461 -411
<< nsubstratencontact >>
rect 1399 315 1403 319
rect 1423 315 1427 319
rect 1449 315 1453 319
rect 1477 315 1481 319
rect 1509 315 1513 319
rect 1107 224 1111 228
rect 1124 224 1128 228
rect 1143 224 1147 228
rect 1175 224 1179 228
rect 1201 224 1205 228
rect 1250 224 1254 228
rect 1282 224 1286 228
rect 775 216 779 220
rect 792 216 796 220
rect 811 216 815 220
rect 843 216 847 220
rect 873 216 877 220
rect 907 216 911 220
rect 939 216 943 220
rect 430 203 434 207
rect 447 203 451 207
rect 466 203 470 207
rect 498 203 502 207
rect 524 203 528 207
rect 543 203 547 207
rect 575 203 579 207
rect 84 160 88 164
rect 101 160 105 164
rect 120 160 124 164
rect 152 160 156 164
rect 1480 151 1484 155
rect 1529 151 1533 155
rect 1561 151 1565 155
rect 1153 81 1157 85
rect 1172 81 1176 85
rect 809 73 813 77
rect 828 73 832 77
rect 105 65 109 69
rect 124 65 128 69
rect 451 68 455 72
rect 470 68 474 72
rect 38 26 42 30
rect 57 26 61 30
rect 173 30 177 34
rect 192 30 196 34
rect 384 29 388 33
rect 403 29 407 33
rect 519 33 523 37
rect 538 33 542 37
rect 742 34 746 38
rect 761 34 765 38
rect 1086 42 1090 46
rect 1105 42 1109 46
rect 1221 46 1225 50
rect 1240 46 1244 50
rect 877 38 881 42
rect 896 38 900 42
rect 255 21 259 25
rect 105 -18 109 -14
rect 124 -18 128 -14
rect 601 24 605 28
rect 451 -15 455 -11
rect 470 -15 474 -11
rect 959 29 963 33
rect 809 -10 813 -6
rect 828 -10 832 -6
rect 1303 37 1307 41
rect 1153 -2 1157 2
rect 1172 -2 1176 2
rect 92 -120 96 -116
rect 109 -120 113 -116
rect 128 -120 132 -116
rect 160 -120 164 -116
rect 747 -149 751 -145
rect 764 -149 768 -145
rect 783 -149 787 -145
rect 815 -149 819 -145
rect 845 -149 849 -145
rect 879 -149 883 -145
rect 911 -149 915 -145
rect 1093 -147 1097 -143
rect 1110 -147 1114 -143
rect 1129 -147 1133 -143
rect 1161 -147 1165 -143
rect 1187 -147 1191 -143
rect 1236 -147 1240 -143
rect 1268 -147 1272 -143
rect 422 -164 426 -160
rect 439 -164 443 -160
rect 458 -164 462 -160
rect 490 -164 494 -160
rect 516 -164 520 -160
rect 535 -164 539 -160
rect 567 -164 571 -160
rect 1346 -348 1350 -344
rect 1370 -348 1374 -344
rect 1396 -348 1400 -344
rect 1424 -348 1428 -344
rect 1456 -348 1460 -344
<< labels >>
rlabel metal1 1462 -379 1462 -379 1 GB
rlabel metal1 1515 284 1515 284 1 GA
rlabel metal1 1568 119 1568 119 7 E
rlabel metal1 -28 367 -28 367 4 a3
rlabel metal1 -11 369 -11 369 5 b3
rlabel metal1 318 367 318 367 5 a2
rlabel metal1 335 367 335 367 5 b2
rlabel metal1 676 367 676 367 5 a1
rlabel metal1 693 366 693 366 1 b1
rlabel metal1 1020 366 1020 366 1 a0
rlabel metal1 1038 366 1038 366 1 b0
rlabel metal1 1441 404 1441 404 5 Vdd
rlabel metal1 1387 -449 1387 -449 1 gnd
<< end >>
