magic
tech scmos
timestamp 1701187352
<< nwell >>
rect 135 109 203 121
rect -70 33 -45 45
rect 137 33 205 45
rect -70 -51 -45 -39
rect 139 -43 207 -31
rect 141 -119 209 -107
<< polysilicon >>
rect 147 119 150 123
rect 162 119 165 123
rect 189 119 191 123
rect 38 92 140 96
rect -59 43 -57 47
rect -59 3 -57 35
rect -59 -7 -57 -5
rect 38 -18 42 92
rect 147 88 150 111
rect 162 96 165 111
rect 161 92 165 96
rect 46 84 133 88
rect 146 84 150 88
rect -59 -41 -57 -37
rect -59 -81 -57 -49
rect -59 -91 -57 -89
rect 46 -99 50 84
rect 147 79 150 84
rect 162 79 165 92
rect 189 79 191 111
rect 147 69 150 71
rect 162 69 165 71
rect 189 69 191 71
rect 149 43 152 47
rect 164 43 167 47
rect 191 43 193 47
rect 69 18 91 22
rect 87 -48 91 18
rect 149 12 152 35
rect 164 20 167 35
rect 163 16 167 20
rect 148 8 152 12
rect 149 3 152 8
rect 164 3 167 16
rect 191 3 193 35
rect 149 -7 152 -5
rect 164 -7 167 -5
rect 191 -7 193 -5
rect 151 -33 154 -29
rect 166 -33 169 -29
rect 193 -33 195 -29
rect 71 -52 137 -48
rect 62 -138 66 -68
rect 71 -132 75 -52
rect 151 -64 154 -41
rect 166 -56 169 -41
rect 165 -60 169 -56
rect 150 -68 154 -64
rect 151 -73 154 -68
rect 166 -73 169 -60
rect 193 -73 195 -41
rect 151 -83 154 -81
rect 166 -83 169 -81
rect 193 -83 195 -81
rect 153 -109 156 -105
rect 168 -109 171 -105
rect 195 -109 197 -105
rect 71 -136 146 -132
rect 153 -140 156 -117
rect 168 -132 171 -117
rect 167 -136 171 -132
rect 152 -144 156 -140
rect 153 -149 156 -144
rect 168 -149 171 -136
rect 195 -149 197 -117
rect 153 -159 156 -157
rect 168 -159 171 -157
rect 195 -159 197 -157
<< ndiffusion >>
rect -69 1 -59 3
rect -69 -3 -67 1
rect -63 -3 -59 1
rect -69 -5 -59 -3
rect -57 1 -47 3
rect -57 -3 -53 1
rect -49 -3 -47 1
rect -57 -5 -47 -3
rect -69 -83 -59 -81
rect -69 -87 -67 -83
rect -63 -87 -59 -83
rect -69 -89 -59 -87
rect -57 -83 -47 -81
rect -57 -87 -53 -83
rect -49 -87 -47 -83
rect -57 -89 -47 -87
rect 137 77 147 79
rect 137 73 139 77
rect 143 73 147 77
rect 137 71 147 73
rect 150 71 162 79
rect 165 77 175 79
rect 165 73 169 77
rect 173 73 175 77
rect 165 71 175 73
rect 179 77 189 79
rect 179 73 181 77
rect 185 73 189 77
rect 179 71 189 73
rect 191 77 201 79
rect 191 73 195 77
rect 199 73 201 77
rect 191 71 201 73
rect 139 1 149 3
rect 139 -3 141 1
rect 145 -3 149 1
rect 139 -5 149 -3
rect 152 -5 164 3
rect 167 1 177 3
rect 167 -3 171 1
rect 175 -3 177 1
rect 167 -5 177 -3
rect 181 1 191 3
rect 181 -3 183 1
rect 187 -3 191 1
rect 181 -5 191 -3
rect 193 1 203 3
rect 193 -3 197 1
rect 201 -3 203 1
rect 193 -5 203 -3
rect 141 -75 151 -73
rect 141 -79 143 -75
rect 147 -79 151 -75
rect 141 -81 151 -79
rect 154 -81 166 -73
rect 169 -75 179 -73
rect 169 -79 173 -75
rect 177 -79 179 -75
rect 169 -81 179 -79
rect 183 -75 193 -73
rect 183 -79 185 -75
rect 189 -79 193 -75
rect 183 -81 193 -79
rect 195 -75 205 -73
rect 195 -79 199 -75
rect 203 -79 205 -75
rect 195 -81 205 -79
rect 143 -151 153 -149
rect 143 -155 145 -151
rect 149 -155 153 -151
rect 143 -157 153 -155
rect 156 -157 168 -149
rect 171 -151 181 -149
rect 171 -155 175 -151
rect 179 -155 181 -151
rect 171 -157 181 -155
rect 185 -151 195 -149
rect 185 -155 187 -151
rect 191 -155 195 -151
rect 185 -157 195 -155
rect 197 -151 207 -149
rect 197 -155 201 -151
rect 205 -155 207 -151
rect 197 -157 207 -155
<< pdiffusion >>
rect 137 117 147 119
rect 137 113 139 117
rect 143 113 147 117
rect 137 111 147 113
rect 150 117 162 119
rect 150 113 154 117
rect 158 113 162 117
rect 150 111 162 113
rect 165 117 175 119
rect 165 113 169 117
rect 173 113 175 117
rect 165 111 175 113
rect 179 117 189 119
rect 179 113 181 117
rect 185 113 189 117
rect 179 111 189 113
rect 191 117 201 119
rect 191 113 195 117
rect 199 113 201 117
rect 191 111 201 113
rect -69 41 -59 43
rect -69 37 -67 41
rect -63 37 -59 41
rect -69 35 -59 37
rect -57 41 -47 43
rect -57 37 -53 41
rect -49 37 -47 41
rect -57 35 -47 37
rect -69 -43 -59 -41
rect -69 -47 -67 -43
rect -63 -47 -59 -43
rect -69 -49 -59 -47
rect -57 -43 -47 -41
rect -57 -47 -53 -43
rect -49 -47 -47 -43
rect -57 -49 -47 -47
rect 139 41 149 43
rect 139 37 141 41
rect 145 37 149 41
rect 139 35 149 37
rect 152 41 164 43
rect 152 37 156 41
rect 160 37 164 41
rect 152 35 164 37
rect 167 41 177 43
rect 167 37 171 41
rect 175 37 177 41
rect 167 35 177 37
rect 181 41 191 43
rect 181 37 183 41
rect 187 37 191 41
rect 181 35 191 37
rect 193 41 203 43
rect 193 37 197 41
rect 201 37 203 41
rect 193 35 203 37
rect 141 -35 151 -33
rect 141 -39 143 -35
rect 147 -39 151 -35
rect 141 -41 151 -39
rect 154 -35 166 -33
rect 154 -39 158 -35
rect 162 -39 166 -35
rect 154 -41 166 -39
rect 169 -35 179 -33
rect 169 -39 173 -35
rect 177 -39 179 -35
rect 169 -41 179 -39
rect 183 -35 193 -33
rect 183 -39 185 -35
rect 189 -39 193 -35
rect 183 -41 193 -39
rect 195 -35 205 -33
rect 195 -39 199 -35
rect 203 -39 205 -35
rect 195 -41 205 -39
rect 143 -111 153 -109
rect 143 -115 145 -111
rect 149 -115 153 -111
rect 143 -117 153 -115
rect 156 -111 168 -109
rect 156 -115 160 -111
rect 164 -115 168 -111
rect 156 -117 168 -115
rect 171 -111 181 -109
rect 171 -115 175 -111
rect 179 -115 181 -111
rect 171 -117 181 -115
rect 185 -111 195 -109
rect 185 -115 187 -111
rect 191 -115 195 -111
rect 185 -117 195 -115
rect 197 -111 207 -109
rect 197 -115 201 -111
rect 205 -115 207 -111
rect 197 -117 207 -115
<< metal1 >>
rect -127 143 236 145
rect -127 141 -41 143
rect -37 141 115 143
rect 119 141 236 143
rect 137 127 144 131
rect 148 127 163 131
rect 167 127 181 131
rect 185 127 195 131
rect 199 127 203 131
rect 139 117 143 127
rect 169 117 173 127
rect 181 117 185 127
rect 154 104 158 113
rect 154 100 173 104
rect 169 96 173 100
rect 195 98 199 113
rect 144 92 157 96
rect 169 92 185 96
rect 195 94 236 98
rect 137 84 142 88
rect 169 77 173 92
rect 195 77 199 94
rect 139 65 143 73
rect 181 65 185 73
rect 137 61 144 65
rect 148 61 165 65
rect 169 61 181 65
rect 185 61 196 65
rect 200 61 201 65
rect -70 51 -67 55
rect -63 51 -53 55
rect -49 51 -47 55
rect 139 51 146 55
rect 150 51 165 55
rect 169 51 183 55
rect 187 51 197 55
rect 201 51 205 55
rect -67 41 -63 51
rect 141 41 145 51
rect 171 41 175 51
rect 183 41 187 51
rect -53 22 -49 37
rect 156 28 160 37
rect 156 24 175 28
rect -127 16 -63 20
rect -53 18 65 22
rect 171 20 175 24
rect 197 22 201 37
rect -87 -20 -83 16
rect -53 1 -49 18
rect 98 16 159 20
rect 171 16 187 20
rect 197 18 236 22
rect 98 -3 102 16
rect -67 -11 -63 -3
rect 60 -7 102 -3
rect 129 8 144 12
rect -68 -15 -67 -11
rect -63 -15 -52 -11
rect -48 -15 -45 -11
rect -87 -22 38 -20
rect 60 -20 64 -7
rect 42 -22 64 -20
rect -87 -24 64 -22
rect -70 -33 -67 -29
rect -63 -33 -53 -29
rect -49 -33 -47 -29
rect -67 -43 -63 -33
rect 129 -35 133 8
rect 171 1 175 16
rect 197 1 201 18
rect 141 -11 145 -3
rect 183 -11 187 -3
rect 139 -15 146 -11
rect 150 -15 167 -11
rect 171 -15 183 -11
rect 187 -15 198 -11
rect 202 -15 203 -11
rect 141 -25 148 -21
rect 152 -25 167 -21
rect 171 -25 185 -21
rect 189 -25 199 -21
rect 203 -25 207 -21
rect 62 -39 133 -35
rect 143 -35 147 -25
rect 173 -35 177 -25
rect 185 -35 189 -25
rect -53 -62 -49 -47
rect 62 -62 66 -39
rect 158 -48 162 -39
rect 141 -52 150 -48
rect 158 -52 177 -48
rect 146 -56 150 -52
rect 173 -56 177 -52
rect 199 -54 203 -39
rect 146 -60 161 -56
rect 173 -60 189 -56
rect 199 -58 236 -54
rect -53 -64 66 -62
rect -127 -68 -63 -64
rect -53 -66 62 -64
rect -87 -103 -83 -68
rect -53 -83 -49 -66
rect 79 -68 146 -64
rect -67 -95 -63 -87
rect -68 -99 -67 -95
rect -63 -99 -52 -95
rect -48 -99 -45 -95
rect 79 -103 83 -68
rect 173 -75 177 -60
rect 199 -75 203 -58
rect 143 -87 147 -79
rect 185 -87 189 -79
rect 141 -91 148 -87
rect 152 -91 169 -87
rect 173 -91 185 -87
rect 189 -91 200 -87
rect 204 -91 205 -87
rect 143 -101 150 -97
rect 154 -101 169 -97
rect 173 -101 187 -97
rect 191 -101 201 -97
rect 205 -101 207 -97
rect -87 -107 83 -103
rect 145 -111 149 -101
rect 175 -111 179 -101
rect 187 -111 191 -101
rect 160 -124 164 -115
rect 160 -128 179 -124
rect 175 -132 179 -128
rect 201 -130 205 -115
rect 150 -136 163 -132
rect 175 -136 191 -132
rect 201 -134 236 -130
rect 66 -142 148 -140
rect 62 -144 148 -142
rect 175 -151 179 -136
rect 201 -151 205 -134
rect 145 -163 149 -155
rect 187 -163 191 -155
rect 143 -167 150 -163
rect 154 -167 171 -163
rect 175 -167 187 -163
rect 191 -167 202 -163
rect 206 -167 207 -163
rect -127 -176 -78 -174
rect -74 -176 220 -174
rect 224 -176 236 -174
rect -127 -178 236 -176
<< metal2 >>
rect -41 55 -37 139
rect -43 51 -37 55
rect -78 -15 -72 -11
rect -78 -95 -74 -15
rect -41 -29 -37 51
rect -43 -33 -37 -29
rect 115 131 119 139
rect 115 127 133 131
rect 115 55 119 127
rect 205 61 224 65
rect 115 51 135 55
rect 115 -21 119 51
rect 220 -11 224 61
rect 207 -15 224 -11
rect 115 -25 137 -21
rect -78 -99 -72 -95
rect 115 -97 119 -25
rect 220 -87 224 -15
rect 209 -91 224 -87
rect -78 -172 -74 -99
rect 115 -101 139 -97
rect 220 -163 224 -91
rect 211 -167 224 -163
rect 220 -172 224 -167
<< ntransistor >>
rect -59 -5 -57 3
rect -59 -89 -57 -81
rect 147 71 150 79
rect 162 71 165 79
rect 189 71 191 79
rect 149 -5 152 3
rect 164 -5 167 3
rect 191 -5 193 3
rect 151 -81 154 -73
rect 166 -81 169 -73
rect 193 -81 195 -73
rect 153 -157 156 -149
rect 168 -157 171 -149
rect 195 -157 197 -149
<< ptransistor >>
rect 147 111 150 119
rect 162 111 165 119
rect 189 111 191 119
rect -59 35 -57 43
rect -59 -49 -57 -41
rect 149 35 152 43
rect 164 35 167 43
rect 191 35 193 43
rect 151 -41 154 -33
rect 166 -41 169 -33
rect 193 -41 195 -33
rect 153 -117 156 -109
rect 168 -117 171 -109
rect 195 -117 197 -109
<< polycontact >>
rect 140 92 144 96
rect -63 16 -59 20
rect 157 92 161 96
rect 185 92 189 96
rect 38 -22 42 -18
rect 133 84 137 88
rect 142 84 146 88
rect -63 -68 -59 -64
rect 65 18 69 22
rect 159 16 163 20
rect 187 16 191 20
rect 144 8 148 12
rect 137 -52 141 -48
rect 46 -103 50 -99
rect 62 -68 66 -64
rect 161 -60 165 -56
rect 189 -60 193 -56
rect 146 -68 150 -64
rect 146 -136 150 -132
rect 62 -142 66 -138
rect 163 -136 167 -132
rect 191 -136 195 -132
rect 148 -144 152 -140
<< ndcontact >>
rect -67 -3 -63 1
rect -53 -3 -49 1
rect -67 -87 -63 -83
rect -53 -87 -49 -83
rect 139 73 143 77
rect 169 73 173 77
rect 181 73 185 77
rect 195 73 199 77
rect 141 -3 145 1
rect 171 -3 175 1
rect 183 -3 187 1
rect 197 -3 201 1
rect 143 -79 147 -75
rect 173 -79 177 -75
rect 185 -79 189 -75
rect 199 -79 203 -75
rect 145 -155 149 -151
rect 175 -155 179 -151
rect 187 -155 191 -151
rect 201 -155 205 -151
<< pdcontact >>
rect 139 113 143 117
rect 154 113 158 117
rect 169 113 173 117
rect 181 113 185 117
rect 195 113 199 117
rect -67 37 -63 41
rect -53 37 -49 41
rect -67 -47 -63 -43
rect -53 -47 -49 -43
rect 141 37 145 41
rect 156 37 160 41
rect 171 37 175 41
rect 183 37 187 41
rect 197 37 201 41
rect 143 -39 147 -35
rect 158 -39 162 -35
rect 173 -39 177 -35
rect 185 -39 189 -35
rect 199 -39 203 -35
rect 145 -115 149 -111
rect 160 -115 164 -111
rect 175 -115 179 -111
rect 187 -115 191 -111
rect 201 -115 205 -111
<< nbccdiffcontact >>
rect 181 127 185 131
rect -67 51 -63 55
rect -67 -33 -63 -29
rect 183 51 187 55
rect 185 -25 189 -21
rect 187 -101 191 -97
<< m2contact >>
rect -41 139 -37 143
rect 115 139 119 143
rect 133 127 137 131
rect 201 61 205 65
rect -47 51 -43 55
rect 135 51 139 55
rect -72 -15 -68 -11
rect -47 -33 -43 -29
rect 203 -15 207 -11
rect 137 -25 141 -21
rect -72 -99 -68 -95
rect 205 -91 209 -87
rect 139 -101 143 -97
rect 207 -167 211 -163
rect -78 -176 -74 -172
rect 220 -176 224 -172
<< psubstratepcontact >>
rect -67 -15 -63 -11
rect -52 -15 -48 -11
rect -67 -99 -63 -95
rect -52 -99 -48 -95
rect 144 61 148 65
rect 165 61 169 65
rect 181 61 185 65
rect 196 61 200 65
rect 146 -15 150 -11
rect 167 -15 171 -11
rect 183 -15 187 -11
rect 198 -15 202 -11
rect 148 -91 152 -87
rect 169 -91 173 -87
rect 185 -91 189 -87
rect 200 -91 204 -87
rect 150 -167 154 -163
rect 171 -167 175 -163
rect 187 -167 191 -163
rect 202 -167 206 -163
<< nsubstratencontact >>
rect 144 127 148 131
rect 163 127 167 131
rect 195 127 199 131
rect -53 51 -49 55
rect -53 -33 -49 -29
rect 146 51 150 55
rect 165 51 169 55
rect 197 51 201 55
rect 148 -25 152 -21
rect 167 -25 171 -21
rect 199 -25 203 -21
rect 150 -101 154 -97
rect 169 -101 173 -97
rect 201 -101 205 -97
<< end >>
