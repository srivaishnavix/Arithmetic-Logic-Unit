* SPICE3 file created from 5ANDGAT.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'


.option scale=1u

M1000 a_2_51# Va Vdd w_n13_49# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1001 a_2_3# Va gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1002 a_17_3# Vb a_2_3# Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=48p ps=20u
M1003 a_2_51# Vd a_2_51# w_n13_49# CMOSP w=8 l=3
+  ad=48p pd=20u as=0.384n ps=0.16m
M1004 Vdd Ve a_2_51# w_n13_49# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1005 Vout a_2_51# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1006 a_2_51# Ve a_47_3# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1007 a_32_3# Vc a_17_3# Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=48p ps=20u
M1008 a_2_51# Vb a_2_51# w_n13_49# CMOSP w=8 l=3
+  ad=48p pd=20u as=0 ps=0
M1009 a_2_51# Vc a_2_51# w_n13_49# CMOSP w=8 l=3
+  ad=48p pd=20u as=0 ps=0
M1010 Vout a_2_51# Vdd w_n13_49# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1011 a_47_3# Vd a_32_3# Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=48p ps=20u
C0 gnd 0 20.116001f 
C1 Vout 0 7.895999f 
C2 a_2_51# 0 32.975998f 
C3 Ve 0 25.882f 
C4 Vd 0 23.626f 
C5 Vc 0 21.369999f 
C6 Vb 0 19.114f 
C7 Va 0 16.858f 
C8 Vdd 0 21.619999f 


Va Va gnd 1
Vb Vb gnd 1
Vc Vc gnd 1
Vd Vd gnd 0
Ve Ve gnd 1


.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(Va) v(Vb)+2 v(Vc)+4 v(Vd)+6 v(Ve)+8 v(Vout)+10 
.end
.endc