magic
tech scmos
timestamp 1701015884
<< nwell >>
rect -22 56 20 68
rect 213 56 255 68
rect -89 17 -47 29
rect 46 21 88 33
rect 146 17 188 29
rect 281 21 323 33
rect -22 -27 20 -15
rect 213 -27 255 -15
rect -108 -117 -40 -105
rect 144 -117 212 -105
rect 261 -117 329 -105
<< polysilicon >>
rect -144 -2 -140 89
rect -136 6 -132 89
rect -10 66 -7 70
rect 5 66 8 70
rect 225 66 228 70
rect 240 66 243 70
rect -10 35 -7 58
rect 5 43 8 58
rect 4 39 8 43
rect -11 31 -7 35
rect -77 27 -74 31
rect -62 27 -59 31
rect -10 26 -7 31
rect 5 26 8 39
rect 225 35 228 58
rect 240 43 243 58
rect 239 39 243 43
rect 58 31 61 35
rect 73 31 76 35
rect 224 31 228 35
rect -118 10 -107 13
rect -118 -101 -115 10
rect -110 7 -107 10
rect -110 6 -106 7
rect -77 -4 -74 19
rect -62 4 -59 19
rect 158 27 161 31
rect 173 27 176 31
rect -10 16 -7 18
rect 5 16 8 18
rect -63 0 -59 4
rect 58 0 61 23
rect 73 8 76 23
rect 225 26 228 31
rect 240 26 243 39
rect 293 31 296 35
rect 308 31 311 35
rect 72 4 76 8
rect -78 -8 -74 -4
rect -110 -11 -106 -10
rect -110 -53 -107 -11
rect -77 -13 -74 -8
rect -62 -13 -59 0
rect 57 -4 61 0
rect 58 -9 61 -4
rect 73 -9 76 4
rect -10 -17 -7 -13
rect 5 -17 8 -13
rect -77 -23 -74 -21
rect -62 -23 -59 -21
rect 58 -19 61 -17
rect 73 -19 76 -17
rect -10 -48 -7 -25
rect 5 -40 8 -25
rect 4 -44 8 -40
rect -11 -52 -7 -48
rect -110 -56 -85 -53
rect -88 -101 -85 -56
rect -10 -57 -7 -52
rect 5 -57 8 -44
rect -10 -67 -7 -65
rect 5 -67 8 -65
rect -118 -104 -93 -101
rect -88 -104 -78 -101
rect -96 -107 -93 -104
rect -81 -107 -78 -104
rect -54 -107 -52 -103
rect -96 -147 -93 -115
rect -81 -147 -78 -115
rect -54 -147 -52 -115
rect -96 -157 -93 -155
rect -81 -157 -78 -155
rect -54 -157 -52 -155
rect -38 -169 -34 -128
rect 97 -138 101 -89
rect 109 -122 113 2
rect 158 -4 161 19
rect 173 4 176 19
rect 225 16 228 18
rect 240 16 243 18
rect 172 0 176 4
rect 293 0 296 23
rect 308 8 311 23
rect 307 4 311 8
rect 157 -8 161 -4
rect 123 -81 127 -10
rect 158 -13 161 -8
rect 173 -13 176 0
rect 292 -4 296 0
rect 293 -9 296 -4
rect 308 -9 311 4
rect 225 -17 228 -13
rect 240 -17 243 -13
rect 158 -23 161 -21
rect 173 -23 176 -21
rect 293 -19 296 -17
rect 308 -19 311 -17
rect 225 -48 228 -25
rect 240 -40 243 -25
rect 239 -44 243 -40
rect 224 -52 228 -48
rect 225 -57 228 -52
rect 240 -57 243 -44
rect 225 -67 228 -65
rect 240 -67 243 -65
rect 156 -107 159 -103
rect 171 -107 174 -103
rect 198 -107 200 -103
rect 273 -107 276 -103
rect 288 -107 291 -103
rect 315 -107 317 -103
rect 109 -126 111 -122
rect 156 -138 159 -115
rect 171 -130 174 -115
rect 170 -134 174 -130
rect 97 -142 99 -138
rect 155 -142 159 -138
rect 156 -147 159 -142
rect 171 -147 174 -134
rect 198 -147 200 -115
rect 273 -138 276 -115
rect 272 -142 276 -138
rect 273 -147 276 -142
rect 288 -147 291 -115
rect 315 -147 317 -115
rect 156 -157 159 -155
rect 171 -157 174 -155
rect 198 -157 200 -155
rect 273 -157 276 -155
rect 288 -157 291 -155
rect 315 -157 317 -155
rect 273 -159 280 -157
rect 277 -169 280 -159
rect -38 -173 280 -169
rect 350 -180 354 2
<< ndiffusion >>
rect -20 24 -10 26
rect -20 20 -18 24
rect -14 20 -10 24
rect -20 18 -10 20
rect -7 18 5 26
rect 8 24 18 26
rect 8 20 12 24
rect 16 20 18 24
rect 8 18 18 20
rect 215 24 225 26
rect 215 20 217 24
rect 221 20 225 24
rect 48 -11 58 -9
rect -87 -15 -77 -13
rect -87 -19 -85 -15
rect -81 -19 -77 -15
rect -87 -21 -77 -19
rect -74 -21 -62 -13
rect -59 -15 -49 -13
rect -59 -19 -55 -15
rect -51 -19 -49 -15
rect 48 -15 50 -11
rect 54 -15 58 -11
rect 48 -17 58 -15
rect 61 -17 73 -9
rect 76 -11 86 -9
rect 76 -15 80 -11
rect 84 -15 86 -11
rect 76 -17 86 -15
rect -59 -21 -49 -19
rect -20 -59 -10 -57
rect -20 -63 -18 -59
rect -14 -63 -10 -59
rect -20 -65 -10 -63
rect -7 -65 5 -57
rect 8 -59 18 -57
rect 8 -63 12 -59
rect 16 -63 18 -59
rect 8 -65 18 -63
rect -106 -149 -96 -147
rect -106 -153 -104 -149
rect -100 -153 -96 -149
rect -106 -155 -96 -153
rect -93 -155 -81 -147
rect -78 -149 -68 -147
rect -78 -153 -74 -149
rect -70 -153 -68 -149
rect -78 -155 -68 -153
rect -64 -149 -54 -147
rect -64 -153 -62 -149
rect -58 -153 -54 -149
rect -64 -155 -54 -153
rect -52 -149 -42 -147
rect -52 -153 -48 -149
rect -44 -153 -42 -149
rect -52 -155 -42 -153
rect 215 18 225 20
rect 228 18 240 26
rect 243 24 253 26
rect 243 20 247 24
rect 251 20 253 24
rect 243 18 253 20
rect 283 -11 293 -9
rect 148 -15 158 -13
rect 148 -19 150 -15
rect 154 -19 158 -15
rect 148 -21 158 -19
rect 161 -21 173 -13
rect 176 -15 186 -13
rect 176 -19 180 -15
rect 184 -19 186 -15
rect 283 -15 285 -11
rect 289 -15 293 -11
rect 283 -17 293 -15
rect 296 -17 308 -9
rect 311 -11 321 -9
rect 311 -15 315 -11
rect 319 -15 321 -11
rect 311 -17 321 -15
rect 176 -21 186 -19
rect 215 -59 225 -57
rect 215 -63 217 -59
rect 221 -63 225 -59
rect 215 -65 225 -63
rect 228 -65 240 -57
rect 243 -59 253 -57
rect 243 -63 247 -59
rect 251 -63 253 -59
rect 243 -65 253 -63
rect 146 -149 156 -147
rect 146 -153 148 -149
rect 152 -153 156 -149
rect 146 -155 156 -153
rect 159 -155 171 -147
rect 174 -149 184 -147
rect 174 -153 178 -149
rect 182 -153 184 -149
rect 174 -155 184 -153
rect 188 -149 198 -147
rect 188 -153 190 -149
rect 194 -153 198 -149
rect 188 -155 198 -153
rect 200 -149 210 -147
rect 200 -153 204 -149
rect 208 -153 210 -149
rect 200 -155 210 -153
rect 263 -149 273 -147
rect 263 -153 265 -149
rect 269 -153 273 -149
rect 263 -155 273 -153
rect 276 -149 288 -147
rect 276 -153 279 -149
rect 283 -153 288 -149
rect 276 -155 288 -153
rect 291 -149 301 -147
rect 291 -153 295 -149
rect 299 -153 301 -149
rect 291 -155 301 -153
rect 305 -149 315 -147
rect 305 -153 307 -149
rect 311 -153 315 -149
rect 305 -155 315 -153
rect 317 -149 327 -147
rect 317 -153 321 -149
rect 325 -153 327 -149
rect 317 -155 327 -153
<< pdiffusion >>
rect -20 64 -10 66
rect -20 60 -18 64
rect -14 60 -10 64
rect -20 58 -10 60
rect -7 64 5 66
rect -7 60 -3 64
rect 1 60 5 64
rect -7 58 5 60
rect 8 64 18 66
rect 8 60 12 64
rect 16 60 18 64
rect 8 58 18 60
rect 215 64 225 66
rect 215 60 217 64
rect 221 60 225 64
rect 215 58 225 60
rect 228 64 240 66
rect 228 60 232 64
rect 236 60 240 64
rect 228 58 240 60
rect 243 64 253 66
rect 243 60 247 64
rect 251 60 253 64
rect 243 58 253 60
rect -87 25 -77 27
rect -87 21 -85 25
rect -81 21 -77 25
rect -87 19 -77 21
rect -74 25 -62 27
rect -74 21 -70 25
rect -66 21 -62 25
rect -74 19 -62 21
rect -59 25 -49 27
rect 48 29 58 31
rect -59 21 -55 25
rect -51 21 -49 25
rect -59 19 -49 21
rect 48 25 50 29
rect 54 25 58 29
rect 48 23 58 25
rect 61 29 73 31
rect 61 25 65 29
rect 69 25 73 29
rect 61 23 73 25
rect 76 29 86 31
rect 76 25 80 29
rect 84 25 86 29
rect 76 23 86 25
rect 148 25 158 27
rect 148 21 150 25
rect 154 21 158 25
rect 148 19 158 21
rect 161 25 173 27
rect 161 21 165 25
rect 169 21 173 25
rect 161 19 173 21
rect 176 25 186 27
rect 283 29 293 31
rect 176 21 180 25
rect 184 21 186 25
rect 176 19 186 21
rect -20 -19 -10 -17
rect -20 -23 -18 -19
rect -14 -23 -10 -19
rect -20 -25 -10 -23
rect -7 -19 5 -17
rect -7 -23 -3 -19
rect 1 -23 5 -19
rect -7 -25 5 -23
rect 8 -19 18 -17
rect 8 -23 12 -19
rect 16 -23 18 -19
rect 8 -25 18 -23
rect -106 -109 -96 -107
rect -106 -113 -104 -109
rect -100 -113 -96 -109
rect -106 -115 -96 -113
rect -93 -109 -81 -107
rect -93 -113 -89 -109
rect -85 -113 -81 -109
rect -93 -115 -81 -113
rect -78 -109 -68 -107
rect -78 -113 -74 -109
rect -70 -113 -68 -109
rect -78 -115 -68 -113
rect -64 -109 -54 -107
rect -64 -113 -62 -109
rect -58 -113 -54 -109
rect -64 -115 -54 -113
rect -52 -109 -42 -107
rect -52 -113 -48 -109
rect -44 -113 -42 -109
rect -52 -115 -42 -113
rect 283 25 285 29
rect 289 25 293 29
rect 283 23 293 25
rect 296 29 308 31
rect 296 25 300 29
rect 304 25 308 29
rect 296 23 308 25
rect 311 29 321 31
rect 311 25 315 29
rect 319 25 321 29
rect 311 23 321 25
rect 215 -19 225 -17
rect 215 -23 217 -19
rect 221 -23 225 -19
rect 215 -25 225 -23
rect 228 -19 240 -17
rect 228 -23 232 -19
rect 236 -23 240 -19
rect 228 -25 240 -23
rect 243 -19 253 -17
rect 243 -23 247 -19
rect 251 -23 253 -19
rect 243 -25 253 -23
rect 146 -109 156 -107
rect 146 -113 148 -109
rect 152 -113 156 -109
rect 146 -115 156 -113
rect 159 -109 171 -107
rect 159 -113 163 -109
rect 167 -113 171 -109
rect 159 -115 171 -113
rect 174 -109 184 -107
rect 174 -113 178 -109
rect 182 -113 184 -109
rect 174 -115 184 -113
rect 188 -109 198 -107
rect 188 -113 190 -109
rect 194 -113 198 -109
rect 188 -115 198 -113
rect 200 -109 210 -107
rect 200 -113 204 -109
rect 208 -113 210 -109
rect 200 -115 210 -113
rect 263 -109 273 -107
rect 263 -113 265 -109
rect 269 -113 273 -109
rect 263 -115 273 -113
rect 276 -115 288 -107
rect 291 -109 301 -107
rect 291 -113 295 -109
rect 299 -113 301 -109
rect 291 -115 301 -113
rect 305 -109 315 -107
rect 305 -113 307 -109
rect 311 -113 315 -109
rect 305 -115 315 -113
rect 317 -109 327 -107
rect 317 -113 321 -109
rect 325 -113 327 -109
rect 317 -115 327 -113
<< metal1 >>
rect -158 76 -13 78
rect -158 74 -50 76
rect -46 74 -13 76
rect -9 74 6 78
rect 10 76 222 78
rect 10 74 185 76
rect -18 64 -14 74
rect 12 64 16 74
rect -3 51 1 60
rect -3 47 16 51
rect -97 43 -22 47
rect 12 43 16 47
rect 67 43 71 74
rect 189 74 222 76
rect 226 74 241 78
rect 245 76 365 78
rect 245 74 341 76
rect 217 64 221 74
rect 247 64 251 74
rect 232 51 236 60
rect 232 47 251 51
rect 138 43 213 47
rect 247 43 251 47
rect 302 43 306 74
rect 345 74 365 76
rect -132 2 -110 4
rect -97 4 -92 43
rect -26 39 0 43
rect 12 39 32 43
rect 48 39 55 43
rect 59 39 74 43
rect 78 39 88 43
rect -89 35 -80 39
rect -76 35 -61 39
rect -57 35 -52 39
rect -85 25 -81 35
rect -55 25 -51 35
rect -35 31 -15 35
rect -70 12 -66 21
rect -70 8 -51 12
rect -55 4 -51 8
rect -35 4 -31 31
rect 12 24 16 39
rect -18 12 -14 20
rect -20 8 -13 12
rect -9 8 8 12
rect 12 8 16 12
rect 28 8 32 39
rect 50 29 54 39
rect 80 29 84 39
rect 65 16 69 25
rect 65 12 84 16
rect 80 8 84 12
rect 138 8 143 43
rect 209 39 235 43
rect 247 39 267 43
rect 283 39 290 43
rect 294 39 309 43
rect 313 39 323 43
rect 146 35 155 39
rect 159 35 174 39
rect 178 35 183 39
rect 150 25 154 35
rect 180 25 184 35
rect 200 31 220 35
rect 165 12 169 21
rect 165 8 184 12
rect 28 4 68 8
rect 80 6 143 8
rect 80 4 109 6
rect -106 2 -67 4
rect -136 0 -67 2
rect -55 0 -31 4
rect -152 -6 -144 -4
rect -140 -6 -82 -4
rect -152 -8 -110 -6
rect -106 -8 -82 -6
rect -95 -35 -90 -8
rect -55 -15 -51 0
rect -85 -27 -81 -19
rect -87 -31 -80 -27
rect -76 -31 -59 -27
rect -55 -31 -50 -27
rect -95 -39 -40 -35
rect -45 -48 -40 -39
rect -35 -40 -31 0
rect 28 -4 53 0
rect -19 -9 -13 -5
rect -9 -9 6 -5
rect 10 -9 18 -5
rect -18 -19 -14 -9
rect 12 -19 16 -9
rect -3 -32 1 -23
rect -3 -36 16 -32
rect 12 -40 16 -36
rect 28 -40 32 -4
rect 80 -11 84 4
rect 113 4 143 6
rect 180 4 184 8
rect 200 4 204 31
rect 247 24 251 39
rect 217 12 221 20
rect 215 8 222 12
rect 226 8 243 12
rect 247 8 251 12
rect 263 8 267 39
rect 285 29 289 39
rect 315 29 319 39
rect 300 16 304 25
rect 300 12 319 16
rect 315 8 319 12
rect 263 4 303 8
rect 315 6 354 8
rect 315 4 350 6
rect 138 0 168 4
rect 180 0 204 4
rect 123 -6 153 -4
rect 127 -8 153 -6
rect 50 -23 54 -15
rect 50 -27 55 -23
rect 59 -27 76 -23
rect 80 -27 84 -23
rect 140 -35 145 -8
rect 180 -15 184 0
rect 150 -27 154 -19
rect 148 -31 155 -27
rect 159 -31 176 -27
rect 180 -31 185 -27
rect 140 -39 195 -35
rect -35 -44 0 -40
rect 12 -44 32 -40
rect -45 -52 -15 -48
rect 12 -59 16 -44
rect 190 -48 195 -39
rect 200 -40 204 0
rect 263 -4 288 0
rect 216 -9 222 -5
rect 226 -9 241 -5
rect 245 -9 253 -5
rect 217 -19 221 -9
rect 247 -19 251 -9
rect 232 -32 236 -23
rect 232 -36 251 -32
rect 247 -40 251 -36
rect 263 -40 267 -4
rect 315 -11 319 4
rect 285 -23 289 -15
rect 285 -27 290 -23
rect 294 -27 311 -23
rect 315 -27 319 -23
rect 200 -44 235 -40
rect 247 -44 267 -40
rect 190 -52 220 -48
rect 247 -59 251 -44
rect -51 -73 -40 -71
rect -18 -71 -14 -63
rect -36 -73 -13 -71
rect -51 -75 -13 -73
rect -9 -75 8 -71
rect 12 -73 20 -71
rect 24 -73 44 -71
rect 48 -73 195 -71
rect 217 -71 221 -63
rect 199 -73 222 -71
rect 12 -75 222 -73
rect 226 -75 243 -71
rect 247 -73 255 -71
rect 259 -73 279 -71
rect 283 -73 347 -71
rect 247 -75 333 -73
rect 337 -75 347 -73
rect -147 -85 123 -83
rect -147 -87 97 -85
rect -147 -128 -143 -87
rect 101 -87 127 -85
rect -107 -99 -99 -95
rect -95 -99 -80 -95
rect -76 -99 -62 -95
rect -58 -99 -48 -95
rect -44 -99 153 -95
rect 157 -99 172 -95
rect 176 -99 190 -95
rect 194 -99 204 -95
rect 208 -99 270 -95
rect 274 -99 289 -95
rect 293 -99 307 -95
rect 311 -99 321 -95
rect 325 -97 341 -95
rect 345 -97 347 -95
rect 325 -99 347 -97
rect -104 -109 -100 -99
rect -74 -109 -70 -99
rect -62 -109 -58 -99
rect 148 -109 152 -99
rect 178 -109 182 -99
rect 190 -109 194 -99
rect 265 -109 269 -99
rect 307 -109 311 -99
rect -89 -122 -85 -113
rect -89 -126 -70 -122
rect -158 -132 -143 -128
rect -74 -130 -70 -126
rect -48 -128 -44 -113
rect 163 -122 167 -113
rect 204 -122 208 -113
rect 115 -126 155 -122
rect 163 -126 182 -122
rect -74 -134 -58 -130
rect -48 -132 -42 -128
rect 151 -130 155 -126
rect 178 -130 182 -126
rect 204 -126 284 -122
rect -74 -149 -70 -134
rect -48 -149 -44 -132
rect 151 -134 166 -130
rect 178 -134 194 -130
rect 103 -142 151 -138
rect 178 -149 182 -134
rect 204 -149 208 -126
rect 295 -130 299 -113
rect 321 -128 325 -113
rect 279 -134 311 -130
rect 321 -132 365 -128
rect 261 -142 268 -138
rect 279 -149 283 -134
rect 321 -149 325 -132
rect -104 -161 -100 -153
rect -62 -161 -58 -153
rect 148 -161 152 -153
rect 190 -161 194 -153
rect 265 -161 269 -153
rect 295 -161 299 -153
rect 307 -161 311 -153
rect -158 -165 -99 -161
rect -95 -165 -78 -161
rect -74 -165 -62 -161
rect -58 -165 -47 -161
rect -43 -165 153 -161
rect 157 -165 174 -161
rect 178 -165 190 -161
rect 194 -165 205 -161
rect 209 -165 270 -161
rect 274 -165 291 -161
rect 295 -165 307 -161
rect 311 -165 322 -161
rect 326 -163 333 -161
rect 337 -163 365 -161
rect 326 -165 365 -163
<< metal2 >>
rect -50 39 -46 72
rect 185 39 189 72
rect -48 35 -38 39
rect 187 35 197 39
rect -42 -5 -38 35
rect -42 -9 -23 -5
rect -46 -31 -36 -27
rect -40 -69 -36 -31
rect 20 -69 24 12
rect 193 -5 197 35
rect 193 -9 212 -5
rect 44 -27 46 -23
rect 44 -69 48 -27
rect 189 -31 199 -27
rect 195 -69 199 -31
rect 255 -69 259 12
rect 279 -27 281 -23
rect 279 -69 283 -27
rect 333 -159 337 -77
rect 341 -93 345 72
<< ntransistor >>
rect -10 18 -7 26
rect 5 18 8 26
rect -77 -21 -74 -13
rect -62 -21 -59 -13
rect 58 -17 61 -9
rect 73 -17 76 -9
rect -10 -65 -7 -57
rect 5 -65 8 -57
rect -96 -155 -93 -147
rect -81 -155 -78 -147
rect -54 -155 -52 -147
rect 225 18 228 26
rect 240 18 243 26
rect 158 -21 161 -13
rect 173 -21 176 -13
rect 293 -17 296 -9
rect 308 -17 311 -9
rect 225 -65 228 -57
rect 240 -65 243 -57
rect 156 -155 159 -147
rect 171 -155 174 -147
rect 198 -155 200 -147
rect 273 -155 276 -147
rect 288 -155 291 -147
rect 315 -155 317 -147
<< ptransistor >>
rect -10 58 -7 66
rect 5 58 8 66
rect 225 58 228 66
rect 240 58 243 66
rect -77 19 -74 27
rect -62 19 -59 27
rect 58 23 61 31
rect 73 23 76 31
rect 158 19 161 27
rect 173 19 176 27
rect -10 -25 -7 -17
rect 5 -25 8 -17
rect -96 -115 -93 -107
rect -81 -115 -78 -107
rect -54 -115 -52 -107
rect 293 23 296 31
rect 308 23 311 31
rect 225 -25 228 -17
rect 240 -25 243 -17
rect 156 -115 159 -107
rect 171 -115 174 -107
rect 198 -115 200 -107
rect 273 -115 276 -107
rect 288 -115 291 -107
rect 315 -115 317 -107
<< polycontact >>
rect 0 39 4 43
rect -15 31 -11 35
rect 235 39 239 43
rect 220 31 224 35
rect -136 2 -132 6
rect -144 -6 -140 -2
rect -110 2 -106 6
rect -67 0 -63 4
rect 68 4 72 8
rect -110 -10 -106 -6
rect -82 -8 -78 -4
rect 53 -4 57 0
rect 109 2 113 6
rect 0 -44 4 -40
rect -15 -52 -11 -48
rect 97 -89 101 -85
rect -58 -134 -54 -130
rect -42 -132 -38 -128
rect 168 0 172 4
rect 303 4 307 8
rect 123 -10 127 -6
rect 153 -8 157 -4
rect 288 -4 292 0
rect 350 2 354 6
rect 235 -44 239 -40
rect 220 -52 224 -48
rect 123 -85 127 -81
rect 111 -126 115 -122
rect 166 -134 170 -130
rect 194 -134 198 -130
rect 99 -142 103 -138
rect 151 -142 155 -138
rect 284 -126 288 -122
rect 268 -142 272 -138
rect 311 -134 315 -130
<< ndcontact >>
rect -18 20 -14 24
rect 12 20 16 24
rect 217 20 221 24
rect -85 -19 -81 -15
rect -55 -19 -51 -15
rect 50 -15 54 -11
rect 80 -15 84 -11
rect -18 -63 -14 -59
rect 12 -63 16 -59
rect -104 -153 -100 -149
rect -74 -153 -70 -149
rect -62 -153 -58 -149
rect -48 -153 -44 -149
rect 247 20 251 24
rect 150 -19 154 -15
rect 180 -19 184 -15
rect 285 -15 289 -11
rect 315 -15 319 -11
rect 217 -63 221 -59
rect 247 -63 251 -59
rect 148 -153 152 -149
rect 178 -153 182 -149
rect 190 -153 194 -149
rect 204 -153 208 -149
rect 265 -153 269 -149
rect 279 -153 283 -149
rect 295 -153 299 -149
rect 307 -153 311 -149
rect 321 -153 325 -149
<< pdcontact >>
rect -18 60 -14 64
rect -3 60 1 64
rect 12 60 16 64
rect 217 60 221 64
rect 232 60 236 64
rect 247 60 251 64
rect -85 21 -81 25
rect -70 21 -66 25
rect -55 21 -51 25
rect 50 25 54 29
rect 65 25 69 29
rect 80 25 84 29
rect 150 21 154 25
rect 165 21 169 25
rect 180 21 184 25
rect -18 -23 -14 -19
rect -3 -23 1 -19
rect 12 -23 16 -19
rect -104 -113 -100 -109
rect -89 -113 -85 -109
rect -74 -113 -70 -109
rect -62 -113 -58 -109
rect -48 -113 -44 -109
rect 285 25 289 29
rect 300 25 304 29
rect 315 25 319 29
rect 217 -23 221 -19
rect 232 -23 236 -19
rect 247 -23 251 -19
rect 148 -113 152 -109
rect 163 -113 167 -109
rect 178 -113 182 -109
rect 190 -113 194 -109
rect 204 -113 208 -109
rect 265 -113 269 -109
rect 295 -113 299 -109
rect 307 -113 311 -109
rect 321 -113 325 -109
<< nbccdiffcontact >>
rect -62 -99 -58 -95
rect 190 -99 194 -95
rect 307 -99 311 -95
<< m2contact >>
rect -50 72 -46 76
rect 185 72 189 76
rect 341 72 345 76
rect -52 35 -48 39
rect 16 8 20 12
rect 183 35 187 39
rect -50 -31 -46 -27
rect -23 -9 -19 -5
rect 251 8 255 12
rect 46 -27 50 -23
rect 185 -31 189 -27
rect 212 -9 216 -5
rect 281 -27 285 -23
rect -40 -73 -36 -69
rect 20 -73 24 -69
rect 44 -73 48 -69
rect 195 -73 199 -69
rect 255 -73 259 -69
rect 279 -73 283 -69
rect 333 -77 337 -73
rect 341 -97 345 -93
rect 333 -163 337 -159
<< psubstratepcontact >>
rect -13 8 -9 12
rect 8 8 12 12
rect -80 -31 -76 -27
rect -59 -31 -55 -27
rect 55 -27 59 -23
rect 76 -27 80 -23
rect -13 -75 -9 -71
rect 8 -75 12 -71
rect -99 -165 -95 -161
rect -78 -165 -74 -161
rect -62 -165 -58 -161
rect -47 -165 -43 -161
rect 222 8 226 12
rect 243 8 247 12
rect 155 -31 159 -27
rect 176 -31 180 -27
rect 290 -27 294 -23
rect 311 -27 315 -23
rect 222 -75 226 -71
rect 243 -75 247 -71
rect 153 -165 157 -161
rect 174 -165 178 -161
rect 190 -165 194 -161
rect 205 -165 209 -161
rect 270 -165 274 -161
rect 291 -165 295 -161
rect 307 -165 311 -161
rect 322 -165 326 -161
<< nsubstratencontact >>
rect -13 74 -9 78
rect 6 74 10 78
rect 222 74 226 78
rect 241 74 245 78
rect -80 35 -76 39
rect -61 35 -57 39
rect 55 39 59 43
rect 74 39 78 43
rect 155 35 159 39
rect 174 35 178 39
rect 290 39 294 43
rect 309 39 313 43
rect -13 -9 -9 -5
rect 6 -9 10 -5
rect -99 -99 -95 -95
rect -80 -99 -76 -95
rect -48 -99 -44 -95
rect 222 -9 226 -5
rect 241 -9 245 -5
rect 153 -99 157 -95
rect 172 -99 176 -95
rect 204 -99 208 -95
rect 270 -99 274 -95
rect 289 -99 293 -95
rect 321 -99 325 -95
<< labels >>
rlabel metal1 130 -6 130 -6 1 c
<< end >>
