4Sub gate implementation 

.include TSMC_180nm.txt
.include NAND.sub
.include NOT.sub
.include AND.sub
.include OR.sub
.include XOR.sub
.include XNOR.sub
.include FullAdder.sub
.include Adder.sub
.include 4Sub.sub


.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_c c gnd dc 1

V_in_a3 a3 gnd dc 0
V_in_a2 a2 gnd dc 1
V_in_a1 a1 gnd dc 1
V_in_a0 a0 gnd dc 1
V_in_b3 b3 gnd dc 1
V_in_b2 b2 gnd dc 1
V_in_b1 b1 gnd dc 1
V_in_b0 b0 gnd dc 1

X1 a3 a2 a1 a0 b3 b2 b1 b0 c s3 s2 s1 s0 cout node_x gnd 4Sub

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(a0) v(b0)+2 v(s0)+4 v(a1)+6 v(b1)+8 v(s1)+10 v(a2)+12 v(b2)+14 v(s2)+16 v(a3)+18 v(b3)+20 v(s3)+22 v(cout)+24

.end
.endc
