magic
tech scmos
timestamp 1701020182
<< nwell >>
rect -144 431 -102 443
rect 369 431 411 443
rect 875 431 917 443
rect 1399 431 1441 443
rect -211 392 -169 404
rect -76 396 -34 408
rect 302 392 344 404
rect 437 396 479 408
rect 808 392 850 404
rect 943 396 985 408
rect 1332 392 1374 404
rect 1467 396 1509 408
rect -144 348 -102 360
rect 369 348 411 360
rect 875 348 917 360
rect 1399 348 1441 360
rect 123 247 165 259
rect 358 247 400 259
rect 646 247 688 259
rect 881 247 923 259
rect 1169 247 1211 259
rect 1404 247 1446 259
rect 1692 247 1734 259
rect 1927 247 1969 259
rect 56 208 98 220
rect 191 212 233 224
rect 291 208 333 220
rect 426 212 468 224
rect 579 208 621 220
rect 714 212 756 224
rect 814 208 856 220
rect 949 212 991 224
rect 1102 208 1144 220
rect 1237 212 1279 224
rect 1337 208 1379 220
rect 1472 212 1514 224
rect 1625 208 1667 220
rect 1760 212 1802 224
rect 1860 208 1902 220
rect 1995 212 2037 224
rect 123 164 165 176
rect 358 164 400 176
rect 646 164 688 176
rect 881 164 923 176
rect 1169 164 1211 176
rect 1404 164 1446 176
rect 1692 164 1734 176
rect 1927 164 1969 176
rect 37 74 105 86
rect 289 74 357 86
rect 406 74 474 86
rect 560 74 628 86
rect 812 74 880 86
rect 929 74 997 86
rect 1083 74 1151 86
rect 1335 74 1403 86
rect 1452 74 1520 86
rect 1606 74 1674 86
rect 1858 74 1926 86
rect 1975 74 2043 86
<< polysilicon >>
rect -278 379 -274 470
rect -132 441 -129 445
rect -117 441 -114 445
rect -132 410 -129 433
rect -117 418 -114 433
rect -118 414 -114 418
rect -133 406 -129 410
rect -199 402 -196 406
rect -184 402 -181 406
rect -132 401 -129 406
rect -117 401 -114 414
rect -64 406 -61 410
rect -49 406 -46 410
rect -278 375 -232 379
rect -199 371 -196 394
rect -184 379 -181 394
rect -132 391 -129 393
rect -117 391 -114 393
rect -185 375 -181 379
rect -64 375 -61 398
rect -49 383 -46 398
rect -50 379 -46 383
rect -200 367 -196 371
rect -199 362 -196 367
rect -184 362 -181 375
rect -65 371 -61 375
rect -64 366 -61 371
rect -49 366 -46 379
rect -132 358 -129 362
rect -117 358 -114 362
rect -199 352 -196 354
rect -184 352 -181 354
rect -64 356 -61 358
rect -49 356 -46 358
rect -132 327 -129 350
rect -117 335 -114 350
rect -118 331 -114 335
rect -133 323 -129 327
rect -132 318 -129 323
rect -117 318 -114 331
rect -132 308 -129 310
rect -117 308 -114 310
rect 1 189 5 468
rect 9 197 13 377
rect 280 379 283 470
rect 381 441 384 445
rect 396 441 399 445
rect 381 410 384 433
rect 396 418 399 433
rect 395 414 399 418
rect 380 406 384 410
rect 314 402 317 406
rect 329 402 332 406
rect 381 401 384 406
rect 396 401 399 414
rect 449 406 452 410
rect 464 406 467 410
rect 280 375 281 379
rect 314 371 317 394
rect 329 379 332 394
rect 381 391 384 393
rect 396 391 399 393
rect 328 375 332 379
rect 449 375 452 398
rect 464 383 467 398
rect 463 379 467 383
rect 279 367 281 371
rect 313 367 317 371
rect 279 289 283 367
rect 314 362 317 367
rect 329 362 332 375
rect 448 371 452 375
rect 449 366 452 371
rect 464 366 467 379
rect 381 358 384 362
rect 396 358 399 362
rect 314 352 317 354
rect 329 352 332 354
rect 449 356 452 358
rect 464 356 467 358
rect 381 327 384 350
rect 396 335 399 350
rect 395 331 399 335
rect 380 323 384 327
rect 381 318 384 323
rect 396 318 399 331
rect 381 308 384 310
rect 396 308 399 310
rect 135 257 138 261
rect 150 257 153 261
rect 370 257 373 261
rect 385 257 388 261
rect 135 226 138 249
rect 150 234 153 249
rect 149 230 153 234
rect 134 222 138 226
rect 68 218 71 222
rect 83 218 86 222
rect 135 217 138 222
rect 150 217 153 230
rect 370 226 373 249
rect 385 234 388 249
rect 384 230 388 234
rect 203 222 206 226
rect 218 222 221 226
rect 369 222 373 226
rect 27 201 38 204
rect 27 90 30 201
rect 35 198 38 201
rect 35 197 39 198
rect 68 187 71 210
rect 83 195 86 210
rect 303 218 306 222
rect 318 218 321 222
rect 135 207 138 209
rect 150 207 153 209
rect 82 191 86 195
rect 203 191 206 214
rect 218 199 221 214
rect 370 217 373 222
rect 385 217 388 230
rect 438 222 441 226
rect 453 222 456 226
rect 217 195 221 199
rect 67 183 71 187
rect 35 180 39 181
rect 35 138 38 180
rect 68 178 71 183
rect 83 178 86 191
rect 202 187 206 191
rect 203 182 206 187
rect 218 182 221 195
rect 135 174 138 178
rect 150 174 153 178
rect 68 168 71 170
rect 83 168 86 170
rect 203 172 206 174
rect 218 172 221 174
rect 135 143 138 166
rect 150 151 153 166
rect 149 147 153 151
rect 134 139 138 143
rect 35 135 60 138
rect 57 90 60 135
rect 135 134 138 139
rect 150 134 153 147
rect 135 124 138 126
rect 150 124 153 126
rect 27 87 52 90
rect 57 87 67 90
rect 49 84 52 87
rect 64 84 67 87
rect 91 84 93 88
rect 49 44 52 76
rect 64 44 67 76
rect 91 44 93 76
rect 49 34 52 36
rect 64 34 67 36
rect 91 34 93 36
rect 107 22 111 63
rect 242 53 246 102
rect 254 69 258 193
rect 303 187 306 210
rect 318 195 321 210
rect 370 207 373 209
rect 385 207 388 209
rect 317 191 321 195
rect 438 191 441 214
rect 453 199 456 214
rect 452 195 456 199
rect 302 183 306 187
rect 268 110 272 181
rect 303 178 306 183
rect 318 178 321 191
rect 437 187 441 191
rect 438 182 441 187
rect 453 182 456 195
rect 370 174 373 178
rect 385 174 388 178
rect 303 168 306 170
rect 318 168 321 170
rect 438 172 441 174
rect 453 172 456 174
rect 370 143 373 166
rect 385 151 388 166
rect 384 147 388 151
rect 369 139 373 143
rect 370 134 373 139
rect 385 134 388 147
rect 370 124 373 126
rect 385 124 388 126
rect 301 84 304 88
rect 316 84 319 88
rect 343 84 345 88
rect 418 84 421 88
rect 433 84 436 88
rect 460 84 462 88
rect 254 65 256 69
rect 301 53 304 76
rect 316 61 319 76
rect 315 57 319 61
rect 242 49 244 53
rect 300 49 304 53
rect 301 44 304 49
rect 316 44 319 57
rect 343 44 345 76
rect 418 53 421 76
rect 417 49 421 53
rect 418 44 421 49
rect 433 44 436 76
rect 460 44 462 76
rect 301 34 304 36
rect 316 34 319 36
rect 343 34 345 36
rect 418 34 421 36
rect 433 34 436 36
rect 460 34 462 36
rect 418 32 425 34
rect 422 22 425 32
rect 107 18 425 22
rect 495 11 499 193
rect 524 189 528 470
rect 532 197 536 377
rect 785 379 789 470
rect 887 441 890 445
rect 902 441 905 445
rect 887 410 890 433
rect 902 418 905 433
rect 901 414 905 418
rect 886 406 890 410
rect 820 402 823 406
rect 835 402 838 406
rect 887 401 890 406
rect 902 401 905 414
rect 955 406 958 410
rect 970 406 973 410
rect 785 375 787 379
rect 820 371 823 394
rect 835 379 838 394
rect 887 391 890 393
rect 902 391 905 393
rect 834 375 838 379
rect 955 375 958 398
rect 970 383 973 398
rect 969 379 973 383
rect 785 367 787 371
rect 819 367 823 371
rect 785 289 789 367
rect 820 362 823 367
rect 835 362 838 375
rect 954 371 958 375
rect 955 366 958 371
rect 970 366 973 379
rect 887 358 890 362
rect 902 358 905 362
rect 820 352 823 354
rect 835 352 838 354
rect 955 356 958 358
rect 970 356 973 358
rect 887 327 890 350
rect 902 335 905 350
rect 901 331 905 335
rect 886 323 890 327
rect 887 318 890 323
rect 902 318 905 331
rect 887 308 890 310
rect 902 308 905 310
rect 658 257 661 261
rect 673 257 676 261
rect 893 257 896 261
rect 908 257 911 261
rect 658 226 661 249
rect 673 234 676 249
rect 672 230 676 234
rect 657 222 661 226
rect 591 218 594 222
rect 606 218 609 222
rect 658 217 661 222
rect 673 217 676 230
rect 893 226 896 249
rect 908 234 911 249
rect 907 230 911 234
rect 726 222 729 226
rect 741 222 744 226
rect 892 222 896 226
rect 550 201 561 204
rect 550 90 553 201
rect 558 198 561 201
rect 558 197 562 198
rect 591 187 594 210
rect 606 195 609 210
rect 826 218 829 222
rect 841 218 844 222
rect 658 207 661 209
rect 673 207 676 209
rect 605 191 609 195
rect 726 191 729 214
rect 741 199 744 214
rect 893 217 896 222
rect 908 217 911 230
rect 961 222 964 226
rect 976 222 979 226
rect 740 195 744 199
rect 590 183 594 187
rect 558 180 562 181
rect 558 138 561 180
rect 591 178 594 183
rect 606 178 609 191
rect 725 187 729 191
rect 726 182 729 187
rect 741 182 744 195
rect 658 174 661 178
rect 673 174 676 178
rect 591 168 594 170
rect 606 168 609 170
rect 726 172 729 174
rect 741 172 744 174
rect 658 143 661 166
rect 673 151 676 166
rect 672 147 676 151
rect 657 139 661 143
rect 558 135 583 138
rect 580 90 583 135
rect 658 134 661 139
rect 673 134 676 147
rect 658 124 661 126
rect 673 124 676 126
rect 550 87 575 90
rect 580 87 590 90
rect 572 84 575 87
rect 587 84 590 87
rect 614 84 616 88
rect 572 44 575 76
rect 587 44 590 76
rect 614 44 616 76
rect 572 34 575 36
rect 587 34 590 36
rect 614 34 616 36
rect 630 22 634 63
rect 765 53 769 102
rect 777 69 781 193
rect 826 187 829 210
rect 841 195 844 210
rect 893 207 896 209
rect 908 207 911 209
rect 840 191 844 195
rect 961 191 964 214
rect 976 199 979 214
rect 975 195 979 199
rect 825 183 829 187
rect 791 110 795 181
rect 826 178 829 183
rect 841 178 844 191
rect 960 187 964 191
rect 961 182 964 187
rect 976 182 979 195
rect 893 174 896 178
rect 908 174 911 178
rect 826 168 829 170
rect 841 168 844 170
rect 961 172 964 174
rect 976 172 979 174
rect 893 143 896 166
rect 908 151 911 166
rect 907 147 911 151
rect 892 139 896 143
rect 893 134 896 139
rect 908 134 911 147
rect 893 124 896 126
rect 908 124 911 126
rect 824 84 827 88
rect 839 84 842 88
rect 866 84 868 88
rect 941 84 944 88
rect 956 84 959 88
rect 983 84 985 88
rect 777 65 779 69
rect 824 53 827 76
rect 839 61 842 76
rect 838 57 842 61
rect 765 49 767 53
rect 823 49 827 53
rect 824 44 827 49
rect 839 44 842 57
rect 866 44 868 76
rect 941 53 944 76
rect 940 49 944 53
rect 941 44 944 49
rect 956 44 959 76
rect 983 44 985 76
rect 824 34 827 36
rect 839 34 842 36
rect 866 34 868 36
rect 941 34 944 36
rect 956 34 959 36
rect 983 34 985 36
rect 941 32 948 34
rect 945 22 948 32
rect 630 18 948 22
rect 1018 11 1022 193
rect 1047 189 1051 470
rect 1055 197 1059 377
rect 1309 379 1313 470
rect 1411 441 1414 445
rect 1426 441 1429 445
rect 1411 410 1414 433
rect 1426 418 1429 433
rect 1425 414 1429 418
rect 1410 406 1414 410
rect 1344 402 1347 406
rect 1359 402 1362 406
rect 1411 401 1414 406
rect 1426 401 1429 414
rect 1479 406 1482 410
rect 1494 406 1497 410
rect 1309 375 1311 379
rect 1344 371 1347 394
rect 1359 379 1362 394
rect 1411 391 1414 393
rect 1426 391 1429 393
rect 1358 375 1362 379
rect 1479 375 1482 398
rect 1494 383 1497 398
rect 1493 379 1497 383
rect 1309 367 1311 371
rect 1343 367 1347 371
rect 1309 289 1313 367
rect 1344 362 1347 367
rect 1359 362 1362 375
rect 1478 371 1482 375
rect 1479 366 1482 371
rect 1494 366 1497 379
rect 1411 358 1414 362
rect 1426 358 1429 362
rect 1344 352 1347 354
rect 1359 352 1362 354
rect 1479 356 1482 358
rect 1494 356 1497 358
rect 1411 327 1414 350
rect 1426 335 1429 350
rect 1425 331 1429 335
rect 1410 323 1414 327
rect 1411 318 1414 323
rect 1426 318 1429 331
rect 1411 308 1414 310
rect 1426 308 1429 310
rect 1181 257 1184 261
rect 1196 257 1199 261
rect 1416 257 1419 261
rect 1431 257 1434 261
rect 1181 226 1184 249
rect 1196 234 1199 249
rect 1195 230 1199 234
rect 1180 222 1184 226
rect 1114 218 1117 222
rect 1129 218 1132 222
rect 1181 217 1184 222
rect 1196 217 1199 230
rect 1416 226 1419 249
rect 1431 234 1434 249
rect 1430 230 1434 234
rect 1249 222 1252 226
rect 1264 222 1267 226
rect 1415 222 1419 226
rect 1073 201 1084 204
rect 1073 90 1076 201
rect 1081 198 1084 201
rect 1081 197 1085 198
rect 1114 187 1117 210
rect 1129 195 1132 210
rect 1349 218 1352 222
rect 1364 218 1367 222
rect 1181 207 1184 209
rect 1196 207 1199 209
rect 1128 191 1132 195
rect 1249 191 1252 214
rect 1264 199 1267 214
rect 1416 217 1419 222
rect 1431 217 1434 230
rect 1484 222 1487 226
rect 1499 222 1502 226
rect 1263 195 1267 199
rect 1113 183 1117 187
rect 1081 180 1085 181
rect 1081 138 1084 180
rect 1114 178 1117 183
rect 1129 178 1132 191
rect 1248 187 1252 191
rect 1249 182 1252 187
rect 1264 182 1267 195
rect 1181 174 1184 178
rect 1196 174 1199 178
rect 1114 168 1117 170
rect 1129 168 1132 170
rect 1249 172 1252 174
rect 1264 172 1267 174
rect 1181 143 1184 166
rect 1196 151 1199 166
rect 1195 147 1199 151
rect 1180 139 1184 143
rect 1081 135 1106 138
rect 1103 90 1106 135
rect 1181 134 1184 139
rect 1196 134 1199 147
rect 1181 124 1184 126
rect 1196 124 1199 126
rect 1073 87 1098 90
rect 1103 87 1113 90
rect 1095 84 1098 87
rect 1110 84 1113 87
rect 1137 84 1139 88
rect 1095 44 1098 76
rect 1110 44 1113 76
rect 1137 44 1139 76
rect 1095 34 1098 36
rect 1110 34 1113 36
rect 1137 34 1139 36
rect 1153 22 1157 63
rect 1288 53 1292 102
rect 1300 69 1304 193
rect 1349 187 1352 210
rect 1364 195 1367 210
rect 1416 207 1419 209
rect 1431 207 1434 209
rect 1363 191 1367 195
rect 1484 191 1487 214
rect 1499 199 1502 214
rect 1498 195 1502 199
rect 1348 183 1352 187
rect 1314 110 1318 181
rect 1349 178 1352 183
rect 1364 178 1367 191
rect 1483 187 1487 191
rect 1484 182 1487 187
rect 1499 182 1502 195
rect 1416 174 1419 178
rect 1431 174 1434 178
rect 1349 168 1352 170
rect 1364 168 1367 170
rect 1484 172 1487 174
rect 1499 172 1502 174
rect 1416 143 1419 166
rect 1431 151 1434 166
rect 1430 147 1434 151
rect 1415 139 1419 143
rect 1416 134 1419 139
rect 1431 134 1434 147
rect 1416 124 1419 126
rect 1431 124 1434 126
rect 1347 84 1350 88
rect 1362 84 1365 88
rect 1389 84 1391 88
rect 1464 84 1467 88
rect 1479 84 1482 88
rect 1506 84 1508 88
rect 1300 65 1302 69
rect 1347 53 1350 76
rect 1362 61 1365 76
rect 1361 57 1365 61
rect 1288 49 1290 53
rect 1346 49 1350 53
rect 1347 44 1350 49
rect 1362 44 1365 57
rect 1389 44 1391 76
rect 1464 53 1467 76
rect 1463 49 1467 53
rect 1464 44 1467 49
rect 1479 44 1482 76
rect 1506 44 1508 76
rect 1347 34 1350 36
rect 1362 34 1365 36
rect 1389 34 1391 36
rect 1464 34 1467 36
rect 1479 34 1482 36
rect 1506 34 1508 36
rect 1464 32 1471 34
rect 1468 22 1471 32
rect 1153 18 1471 22
rect 1541 11 1545 193
rect 1570 189 1574 470
rect 1578 197 1582 377
rect 1704 257 1707 261
rect 1719 257 1722 261
rect 1939 257 1942 261
rect 1954 257 1957 261
rect 1704 226 1707 249
rect 1719 234 1722 249
rect 1718 230 1722 234
rect 1703 222 1707 226
rect 1637 218 1640 222
rect 1652 218 1655 222
rect 1704 217 1707 222
rect 1719 217 1722 230
rect 1939 226 1942 249
rect 1954 234 1957 249
rect 1953 230 1957 234
rect 1772 222 1775 226
rect 1787 222 1790 226
rect 1938 222 1942 226
rect 1596 201 1607 204
rect 1596 90 1599 201
rect 1604 198 1607 201
rect 1604 197 1608 198
rect 1637 187 1640 210
rect 1652 195 1655 210
rect 1872 218 1875 222
rect 1887 218 1890 222
rect 1704 207 1707 209
rect 1719 207 1722 209
rect 1651 191 1655 195
rect 1772 191 1775 214
rect 1787 199 1790 214
rect 1939 217 1942 222
rect 1954 217 1957 230
rect 2007 222 2010 226
rect 2022 222 2025 226
rect 1786 195 1790 199
rect 1636 183 1640 187
rect 1604 180 1608 181
rect 1604 138 1607 180
rect 1637 178 1640 183
rect 1652 178 1655 191
rect 1771 187 1775 191
rect 1772 182 1775 187
rect 1787 182 1790 195
rect 1704 174 1707 178
rect 1719 174 1722 178
rect 1637 168 1640 170
rect 1652 168 1655 170
rect 1772 172 1775 174
rect 1787 172 1790 174
rect 1704 143 1707 166
rect 1719 151 1722 166
rect 1718 147 1722 151
rect 1703 139 1707 143
rect 1604 135 1629 138
rect 1626 90 1629 135
rect 1704 134 1707 139
rect 1719 134 1722 147
rect 1704 124 1707 126
rect 1719 124 1722 126
rect 1596 87 1621 90
rect 1626 87 1636 90
rect 1618 84 1621 87
rect 1633 84 1636 87
rect 1660 84 1662 88
rect 1618 44 1621 76
rect 1633 44 1636 76
rect 1660 44 1662 76
rect 1618 34 1621 36
rect 1633 34 1636 36
rect 1660 34 1662 36
rect 1676 22 1680 63
rect 1811 53 1815 102
rect 1823 69 1827 193
rect 1872 187 1875 210
rect 1887 195 1890 210
rect 1939 207 1942 209
rect 1954 207 1957 209
rect 1886 191 1890 195
rect 2007 191 2010 214
rect 2022 199 2025 214
rect 2021 195 2025 199
rect 1871 183 1875 187
rect 1837 110 1841 181
rect 1872 178 1875 183
rect 1887 178 1890 191
rect 2006 187 2010 191
rect 2007 182 2010 187
rect 2022 182 2025 195
rect 1939 174 1942 178
rect 1954 174 1957 178
rect 1872 168 1875 170
rect 1887 168 1890 170
rect 2007 172 2010 174
rect 2022 172 2025 174
rect 1939 143 1942 166
rect 1954 151 1957 166
rect 1953 147 1957 151
rect 1938 139 1942 143
rect 1939 134 1942 139
rect 1954 134 1957 147
rect 1939 124 1942 126
rect 1954 124 1957 126
rect 1870 84 1873 88
rect 1885 84 1888 88
rect 1912 84 1914 88
rect 1987 84 1990 88
rect 2002 84 2005 88
rect 2029 84 2031 88
rect 1823 65 1825 69
rect 1870 53 1873 76
rect 1885 61 1888 76
rect 1884 57 1888 61
rect 1811 49 1813 53
rect 1869 49 1873 53
rect 1870 44 1873 49
rect 1885 44 1888 57
rect 1912 44 1914 76
rect 1987 53 1990 76
rect 1986 49 1990 53
rect 1987 44 1990 49
rect 2002 44 2005 76
rect 2029 44 2031 76
rect 1870 34 1873 36
rect 1885 34 1888 36
rect 1912 34 1914 36
rect 1987 34 1990 36
rect 2002 34 2005 36
rect 2029 34 2031 36
rect 1987 32 1994 34
rect 1991 22 1994 32
rect 1676 18 1994 22
rect 2064 11 2068 193
<< ndiffusion >>
rect -142 399 -132 401
rect -142 395 -140 399
rect -136 395 -132 399
rect -142 393 -132 395
rect -129 393 -117 401
rect -114 399 -104 401
rect -114 395 -110 399
rect -106 395 -104 399
rect -114 393 -104 395
rect -74 364 -64 366
rect -209 360 -199 362
rect -209 356 -207 360
rect -203 356 -199 360
rect -209 354 -199 356
rect -196 354 -184 362
rect -181 360 -171 362
rect -181 356 -177 360
rect -173 356 -171 360
rect -74 360 -72 364
rect -68 360 -64 364
rect -74 358 -64 360
rect -61 358 -49 366
rect -46 364 -36 366
rect -46 360 -42 364
rect -38 360 -36 364
rect -46 358 -36 360
rect -181 354 -171 356
rect -142 316 -132 318
rect -142 312 -140 316
rect -136 312 -132 316
rect -142 310 -132 312
rect -129 310 -117 318
rect -114 316 -104 318
rect -114 312 -110 316
rect -106 312 -104 316
rect -114 310 -104 312
rect 371 399 381 401
rect 371 395 373 399
rect 377 395 381 399
rect 371 393 381 395
rect 384 393 396 401
rect 399 399 409 401
rect 399 395 403 399
rect 407 395 409 399
rect 399 393 409 395
rect 439 364 449 366
rect 304 360 314 362
rect 304 356 306 360
rect 310 356 314 360
rect 304 354 314 356
rect 317 354 329 362
rect 332 360 342 362
rect 332 356 336 360
rect 340 356 342 360
rect 439 360 441 364
rect 445 360 449 364
rect 439 358 449 360
rect 452 358 464 366
rect 467 364 477 366
rect 467 360 471 364
rect 475 360 477 364
rect 467 358 477 360
rect 332 354 342 356
rect 371 316 381 318
rect 371 312 373 316
rect 377 312 381 316
rect 371 310 381 312
rect 384 310 396 318
rect 399 316 409 318
rect 399 312 403 316
rect 407 312 409 316
rect 399 310 409 312
rect 125 215 135 217
rect 125 211 127 215
rect 131 211 135 215
rect 125 209 135 211
rect 138 209 150 217
rect 153 215 163 217
rect 153 211 157 215
rect 161 211 163 215
rect 153 209 163 211
rect 360 215 370 217
rect 360 211 362 215
rect 366 211 370 215
rect 193 180 203 182
rect 58 176 68 178
rect 58 172 60 176
rect 64 172 68 176
rect 58 170 68 172
rect 71 170 83 178
rect 86 176 96 178
rect 86 172 90 176
rect 94 172 96 176
rect 193 176 195 180
rect 199 176 203 180
rect 193 174 203 176
rect 206 174 218 182
rect 221 180 231 182
rect 221 176 225 180
rect 229 176 231 180
rect 221 174 231 176
rect 86 170 96 172
rect 125 132 135 134
rect 125 128 127 132
rect 131 128 135 132
rect 125 126 135 128
rect 138 126 150 134
rect 153 132 163 134
rect 153 128 157 132
rect 161 128 163 132
rect 153 126 163 128
rect 39 42 49 44
rect 39 38 41 42
rect 45 38 49 42
rect 39 36 49 38
rect 52 36 64 44
rect 67 42 77 44
rect 67 38 71 42
rect 75 38 77 42
rect 67 36 77 38
rect 81 42 91 44
rect 81 38 83 42
rect 87 38 91 42
rect 81 36 91 38
rect 93 42 103 44
rect 93 38 97 42
rect 101 38 103 42
rect 93 36 103 38
rect 360 209 370 211
rect 373 209 385 217
rect 388 215 398 217
rect 388 211 392 215
rect 396 211 398 215
rect 388 209 398 211
rect 428 180 438 182
rect 293 176 303 178
rect 293 172 295 176
rect 299 172 303 176
rect 293 170 303 172
rect 306 170 318 178
rect 321 176 331 178
rect 321 172 325 176
rect 329 172 331 176
rect 428 176 430 180
rect 434 176 438 180
rect 428 174 438 176
rect 441 174 453 182
rect 456 180 466 182
rect 456 176 460 180
rect 464 176 466 180
rect 456 174 466 176
rect 321 170 331 172
rect 360 132 370 134
rect 360 128 362 132
rect 366 128 370 132
rect 360 126 370 128
rect 373 126 385 134
rect 388 132 398 134
rect 388 128 392 132
rect 396 128 398 132
rect 388 126 398 128
rect 291 42 301 44
rect 291 38 293 42
rect 297 38 301 42
rect 291 36 301 38
rect 304 36 316 44
rect 319 42 329 44
rect 319 38 323 42
rect 327 38 329 42
rect 319 36 329 38
rect 333 42 343 44
rect 333 38 335 42
rect 339 38 343 42
rect 333 36 343 38
rect 345 42 355 44
rect 345 38 349 42
rect 353 38 355 42
rect 345 36 355 38
rect 408 42 418 44
rect 408 38 410 42
rect 414 38 418 42
rect 408 36 418 38
rect 421 42 433 44
rect 421 38 424 42
rect 428 38 433 42
rect 421 36 433 38
rect 436 42 446 44
rect 436 38 440 42
rect 444 38 446 42
rect 436 36 446 38
rect 450 42 460 44
rect 450 38 452 42
rect 456 38 460 42
rect 450 36 460 38
rect 462 42 472 44
rect 462 38 466 42
rect 470 38 472 42
rect 462 36 472 38
rect 877 399 887 401
rect 877 395 879 399
rect 883 395 887 399
rect 877 393 887 395
rect 890 393 902 401
rect 905 399 915 401
rect 905 395 909 399
rect 913 395 915 399
rect 905 393 915 395
rect 945 364 955 366
rect 810 360 820 362
rect 810 356 812 360
rect 816 356 820 360
rect 810 354 820 356
rect 823 354 835 362
rect 838 360 848 362
rect 838 356 842 360
rect 846 356 848 360
rect 945 360 947 364
rect 951 360 955 364
rect 945 358 955 360
rect 958 358 970 366
rect 973 364 983 366
rect 973 360 977 364
rect 981 360 983 364
rect 973 358 983 360
rect 838 354 848 356
rect 877 316 887 318
rect 877 312 879 316
rect 883 312 887 316
rect 877 310 887 312
rect 890 310 902 318
rect 905 316 915 318
rect 905 312 909 316
rect 913 312 915 316
rect 905 310 915 312
rect 648 215 658 217
rect 648 211 650 215
rect 654 211 658 215
rect 648 209 658 211
rect 661 209 673 217
rect 676 215 686 217
rect 676 211 680 215
rect 684 211 686 215
rect 676 209 686 211
rect 883 215 893 217
rect 883 211 885 215
rect 889 211 893 215
rect 716 180 726 182
rect 581 176 591 178
rect 581 172 583 176
rect 587 172 591 176
rect 581 170 591 172
rect 594 170 606 178
rect 609 176 619 178
rect 609 172 613 176
rect 617 172 619 176
rect 716 176 718 180
rect 722 176 726 180
rect 716 174 726 176
rect 729 174 741 182
rect 744 180 754 182
rect 744 176 748 180
rect 752 176 754 180
rect 744 174 754 176
rect 609 170 619 172
rect 648 132 658 134
rect 648 128 650 132
rect 654 128 658 132
rect 648 126 658 128
rect 661 126 673 134
rect 676 132 686 134
rect 676 128 680 132
rect 684 128 686 132
rect 676 126 686 128
rect 562 42 572 44
rect 562 38 564 42
rect 568 38 572 42
rect 562 36 572 38
rect 575 36 587 44
rect 590 42 600 44
rect 590 38 594 42
rect 598 38 600 42
rect 590 36 600 38
rect 604 42 614 44
rect 604 38 606 42
rect 610 38 614 42
rect 604 36 614 38
rect 616 42 626 44
rect 616 38 620 42
rect 624 38 626 42
rect 616 36 626 38
rect 883 209 893 211
rect 896 209 908 217
rect 911 215 921 217
rect 911 211 915 215
rect 919 211 921 215
rect 911 209 921 211
rect 951 180 961 182
rect 816 176 826 178
rect 816 172 818 176
rect 822 172 826 176
rect 816 170 826 172
rect 829 170 841 178
rect 844 176 854 178
rect 844 172 848 176
rect 852 172 854 176
rect 951 176 953 180
rect 957 176 961 180
rect 951 174 961 176
rect 964 174 976 182
rect 979 180 989 182
rect 979 176 983 180
rect 987 176 989 180
rect 979 174 989 176
rect 844 170 854 172
rect 883 132 893 134
rect 883 128 885 132
rect 889 128 893 132
rect 883 126 893 128
rect 896 126 908 134
rect 911 132 921 134
rect 911 128 915 132
rect 919 128 921 132
rect 911 126 921 128
rect 814 42 824 44
rect 814 38 816 42
rect 820 38 824 42
rect 814 36 824 38
rect 827 36 839 44
rect 842 42 852 44
rect 842 38 846 42
rect 850 38 852 42
rect 842 36 852 38
rect 856 42 866 44
rect 856 38 858 42
rect 862 38 866 42
rect 856 36 866 38
rect 868 42 878 44
rect 868 38 872 42
rect 876 38 878 42
rect 868 36 878 38
rect 931 42 941 44
rect 931 38 933 42
rect 937 38 941 42
rect 931 36 941 38
rect 944 42 956 44
rect 944 38 947 42
rect 951 38 956 42
rect 944 36 956 38
rect 959 42 969 44
rect 959 38 963 42
rect 967 38 969 42
rect 959 36 969 38
rect 973 42 983 44
rect 973 38 975 42
rect 979 38 983 42
rect 973 36 983 38
rect 985 42 995 44
rect 985 38 989 42
rect 993 38 995 42
rect 985 36 995 38
rect 1401 399 1411 401
rect 1401 395 1403 399
rect 1407 395 1411 399
rect 1401 393 1411 395
rect 1414 393 1426 401
rect 1429 399 1439 401
rect 1429 395 1433 399
rect 1437 395 1439 399
rect 1429 393 1439 395
rect 1469 364 1479 366
rect 1334 360 1344 362
rect 1334 356 1336 360
rect 1340 356 1344 360
rect 1334 354 1344 356
rect 1347 354 1359 362
rect 1362 360 1372 362
rect 1362 356 1366 360
rect 1370 356 1372 360
rect 1469 360 1471 364
rect 1475 360 1479 364
rect 1469 358 1479 360
rect 1482 358 1494 366
rect 1497 364 1507 366
rect 1497 360 1501 364
rect 1505 360 1507 364
rect 1497 358 1507 360
rect 1362 354 1372 356
rect 1401 316 1411 318
rect 1401 312 1403 316
rect 1407 312 1411 316
rect 1401 310 1411 312
rect 1414 310 1426 318
rect 1429 316 1439 318
rect 1429 312 1433 316
rect 1437 312 1439 316
rect 1429 310 1439 312
rect 1171 215 1181 217
rect 1171 211 1173 215
rect 1177 211 1181 215
rect 1171 209 1181 211
rect 1184 209 1196 217
rect 1199 215 1209 217
rect 1199 211 1203 215
rect 1207 211 1209 215
rect 1199 209 1209 211
rect 1406 215 1416 217
rect 1406 211 1408 215
rect 1412 211 1416 215
rect 1239 180 1249 182
rect 1104 176 1114 178
rect 1104 172 1106 176
rect 1110 172 1114 176
rect 1104 170 1114 172
rect 1117 170 1129 178
rect 1132 176 1142 178
rect 1132 172 1136 176
rect 1140 172 1142 176
rect 1239 176 1241 180
rect 1245 176 1249 180
rect 1239 174 1249 176
rect 1252 174 1264 182
rect 1267 180 1277 182
rect 1267 176 1271 180
rect 1275 176 1277 180
rect 1267 174 1277 176
rect 1132 170 1142 172
rect 1171 132 1181 134
rect 1171 128 1173 132
rect 1177 128 1181 132
rect 1171 126 1181 128
rect 1184 126 1196 134
rect 1199 132 1209 134
rect 1199 128 1203 132
rect 1207 128 1209 132
rect 1199 126 1209 128
rect 1085 42 1095 44
rect 1085 38 1087 42
rect 1091 38 1095 42
rect 1085 36 1095 38
rect 1098 36 1110 44
rect 1113 42 1123 44
rect 1113 38 1117 42
rect 1121 38 1123 42
rect 1113 36 1123 38
rect 1127 42 1137 44
rect 1127 38 1129 42
rect 1133 38 1137 42
rect 1127 36 1137 38
rect 1139 42 1149 44
rect 1139 38 1143 42
rect 1147 38 1149 42
rect 1139 36 1149 38
rect 1406 209 1416 211
rect 1419 209 1431 217
rect 1434 215 1444 217
rect 1434 211 1438 215
rect 1442 211 1444 215
rect 1434 209 1444 211
rect 1474 180 1484 182
rect 1339 176 1349 178
rect 1339 172 1341 176
rect 1345 172 1349 176
rect 1339 170 1349 172
rect 1352 170 1364 178
rect 1367 176 1377 178
rect 1367 172 1371 176
rect 1375 172 1377 176
rect 1474 176 1476 180
rect 1480 176 1484 180
rect 1474 174 1484 176
rect 1487 174 1499 182
rect 1502 180 1512 182
rect 1502 176 1506 180
rect 1510 176 1512 180
rect 1502 174 1512 176
rect 1367 170 1377 172
rect 1406 132 1416 134
rect 1406 128 1408 132
rect 1412 128 1416 132
rect 1406 126 1416 128
rect 1419 126 1431 134
rect 1434 132 1444 134
rect 1434 128 1438 132
rect 1442 128 1444 132
rect 1434 126 1444 128
rect 1337 42 1347 44
rect 1337 38 1339 42
rect 1343 38 1347 42
rect 1337 36 1347 38
rect 1350 36 1362 44
rect 1365 42 1375 44
rect 1365 38 1369 42
rect 1373 38 1375 42
rect 1365 36 1375 38
rect 1379 42 1389 44
rect 1379 38 1381 42
rect 1385 38 1389 42
rect 1379 36 1389 38
rect 1391 42 1401 44
rect 1391 38 1395 42
rect 1399 38 1401 42
rect 1391 36 1401 38
rect 1454 42 1464 44
rect 1454 38 1456 42
rect 1460 38 1464 42
rect 1454 36 1464 38
rect 1467 42 1479 44
rect 1467 38 1470 42
rect 1474 38 1479 42
rect 1467 36 1479 38
rect 1482 42 1492 44
rect 1482 38 1486 42
rect 1490 38 1492 42
rect 1482 36 1492 38
rect 1496 42 1506 44
rect 1496 38 1498 42
rect 1502 38 1506 42
rect 1496 36 1506 38
rect 1508 42 1518 44
rect 1508 38 1512 42
rect 1516 38 1518 42
rect 1508 36 1518 38
rect 1694 215 1704 217
rect 1694 211 1696 215
rect 1700 211 1704 215
rect 1694 209 1704 211
rect 1707 209 1719 217
rect 1722 215 1732 217
rect 1722 211 1726 215
rect 1730 211 1732 215
rect 1722 209 1732 211
rect 1929 215 1939 217
rect 1929 211 1931 215
rect 1935 211 1939 215
rect 1762 180 1772 182
rect 1627 176 1637 178
rect 1627 172 1629 176
rect 1633 172 1637 176
rect 1627 170 1637 172
rect 1640 170 1652 178
rect 1655 176 1665 178
rect 1655 172 1659 176
rect 1663 172 1665 176
rect 1762 176 1764 180
rect 1768 176 1772 180
rect 1762 174 1772 176
rect 1775 174 1787 182
rect 1790 180 1800 182
rect 1790 176 1794 180
rect 1798 176 1800 180
rect 1790 174 1800 176
rect 1655 170 1665 172
rect 1694 132 1704 134
rect 1694 128 1696 132
rect 1700 128 1704 132
rect 1694 126 1704 128
rect 1707 126 1719 134
rect 1722 132 1732 134
rect 1722 128 1726 132
rect 1730 128 1732 132
rect 1722 126 1732 128
rect 1608 42 1618 44
rect 1608 38 1610 42
rect 1614 38 1618 42
rect 1608 36 1618 38
rect 1621 36 1633 44
rect 1636 42 1646 44
rect 1636 38 1640 42
rect 1644 38 1646 42
rect 1636 36 1646 38
rect 1650 42 1660 44
rect 1650 38 1652 42
rect 1656 38 1660 42
rect 1650 36 1660 38
rect 1662 42 1672 44
rect 1662 38 1666 42
rect 1670 38 1672 42
rect 1662 36 1672 38
rect 1929 209 1939 211
rect 1942 209 1954 217
rect 1957 215 1967 217
rect 1957 211 1961 215
rect 1965 211 1967 215
rect 1957 209 1967 211
rect 1997 180 2007 182
rect 1862 176 1872 178
rect 1862 172 1864 176
rect 1868 172 1872 176
rect 1862 170 1872 172
rect 1875 170 1887 178
rect 1890 176 1900 178
rect 1890 172 1894 176
rect 1898 172 1900 176
rect 1997 176 1999 180
rect 2003 176 2007 180
rect 1997 174 2007 176
rect 2010 174 2022 182
rect 2025 180 2035 182
rect 2025 176 2029 180
rect 2033 176 2035 180
rect 2025 174 2035 176
rect 1890 170 1900 172
rect 1929 132 1939 134
rect 1929 128 1931 132
rect 1935 128 1939 132
rect 1929 126 1939 128
rect 1942 126 1954 134
rect 1957 132 1967 134
rect 1957 128 1961 132
rect 1965 128 1967 132
rect 1957 126 1967 128
rect 1860 42 1870 44
rect 1860 38 1862 42
rect 1866 38 1870 42
rect 1860 36 1870 38
rect 1873 36 1885 44
rect 1888 42 1898 44
rect 1888 38 1892 42
rect 1896 38 1898 42
rect 1888 36 1898 38
rect 1902 42 1912 44
rect 1902 38 1904 42
rect 1908 38 1912 42
rect 1902 36 1912 38
rect 1914 42 1924 44
rect 1914 38 1918 42
rect 1922 38 1924 42
rect 1914 36 1924 38
rect 1977 42 1987 44
rect 1977 38 1979 42
rect 1983 38 1987 42
rect 1977 36 1987 38
rect 1990 42 2002 44
rect 1990 38 1993 42
rect 1997 38 2002 42
rect 1990 36 2002 38
rect 2005 42 2015 44
rect 2005 38 2009 42
rect 2013 38 2015 42
rect 2005 36 2015 38
rect 2019 42 2029 44
rect 2019 38 2021 42
rect 2025 38 2029 42
rect 2019 36 2029 38
rect 2031 42 2041 44
rect 2031 38 2035 42
rect 2039 38 2041 42
rect 2031 36 2041 38
<< pdiffusion >>
rect -142 439 -132 441
rect -142 435 -140 439
rect -136 435 -132 439
rect -142 433 -132 435
rect -129 439 -117 441
rect -129 435 -125 439
rect -121 435 -117 439
rect -129 433 -117 435
rect -114 439 -104 441
rect -114 435 -110 439
rect -106 435 -104 439
rect -114 433 -104 435
rect -209 400 -199 402
rect -209 396 -207 400
rect -203 396 -199 400
rect -209 394 -199 396
rect -196 400 -184 402
rect -196 396 -192 400
rect -188 396 -184 400
rect -196 394 -184 396
rect -181 400 -171 402
rect -74 404 -64 406
rect -181 396 -177 400
rect -173 396 -171 400
rect -181 394 -171 396
rect -74 400 -72 404
rect -68 400 -64 404
rect -74 398 -64 400
rect -61 404 -49 406
rect -61 400 -57 404
rect -53 400 -49 404
rect -61 398 -49 400
rect -46 404 -36 406
rect -46 400 -42 404
rect -38 400 -36 404
rect -46 398 -36 400
rect -142 356 -132 358
rect -142 352 -140 356
rect -136 352 -132 356
rect -142 350 -132 352
rect -129 356 -117 358
rect -129 352 -125 356
rect -121 352 -117 356
rect -129 350 -117 352
rect -114 356 -104 358
rect -114 352 -110 356
rect -106 352 -104 356
rect -114 350 -104 352
rect 371 439 381 441
rect 371 435 373 439
rect 377 435 381 439
rect 371 433 381 435
rect 384 439 396 441
rect 384 435 388 439
rect 392 435 396 439
rect 384 433 396 435
rect 399 439 409 441
rect 399 435 403 439
rect 407 435 409 439
rect 399 433 409 435
rect 304 400 314 402
rect 304 396 306 400
rect 310 396 314 400
rect 304 394 314 396
rect 317 400 329 402
rect 317 396 321 400
rect 325 396 329 400
rect 317 394 329 396
rect 332 400 342 402
rect 439 404 449 406
rect 332 396 336 400
rect 340 396 342 400
rect 332 394 342 396
rect 439 400 441 404
rect 445 400 449 404
rect 439 398 449 400
rect 452 404 464 406
rect 452 400 456 404
rect 460 400 464 404
rect 452 398 464 400
rect 467 404 477 406
rect 467 400 471 404
rect 475 400 477 404
rect 467 398 477 400
rect 371 356 381 358
rect 371 352 373 356
rect 377 352 381 356
rect 371 350 381 352
rect 384 356 396 358
rect 384 352 388 356
rect 392 352 396 356
rect 384 350 396 352
rect 399 356 409 358
rect 399 352 403 356
rect 407 352 409 356
rect 399 350 409 352
rect 125 255 135 257
rect 125 251 127 255
rect 131 251 135 255
rect 125 249 135 251
rect 138 255 150 257
rect 138 251 142 255
rect 146 251 150 255
rect 138 249 150 251
rect 153 255 163 257
rect 153 251 157 255
rect 161 251 163 255
rect 153 249 163 251
rect 360 255 370 257
rect 360 251 362 255
rect 366 251 370 255
rect 360 249 370 251
rect 373 255 385 257
rect 373 251 377 255
rect 381 251 385 255
rect 373 249 385 251
rect 388 255 398 257
rect 388 251 392 255
rect 396 251 398 255
rect 388 249 398 251
rect 58 216 68 218
rect 58 212 60 216
rect 64 212 68 216
rect 58 210 68 212
rect 71 216 83 218
rect 71 212 75 216
rect 79 212 83 216
rect 71 210 83 212
rect 86 216 96 218
rect 193 220 203 222
rect 86 212 90 216
rect 94 212 96 216
rect 86 210 96 212
rect 193 216 195 220
rect 199 216 203 220
rect 193 214 203 216
rect 206 220 218 222
rect 206 216 210 220
rect 214 216 218 220
rect 206 214 218 216
rect 221 220 231 222
rect 221 216 225 220
rect 229 216 231 220
rect 221 214 231 216
rect 293 216 303 218
rect 293 212 295 216
rect 299 212 303 216
rect 293 210 303 212
rect 306 216 318 218
rect 306 212 310 216
rect 314 212 318 216
rect 306 210 318 212
rect 321 216 331 218
rect 428 220 438 222
rect 321 212 325 216
rect 329 212 331 216
rect 321 210 331 212
rect 125 172 135 174
rect 125 168 127 172
rect 131 168 135 172
rect 125 166 135 168
rect 138 172 150 174
rect 138 168 142 172
rect 146 168 150 172
rect 138 166 150 168
rect 153 172 163 174
rect 153 168 157 172
rect 161 168 163 172
rect 153 166 163 168
rect 39 82 49 84
rect 39 78 41 82
rect 45 78 49 82
rect 39 76 49 78
rect 52 82 64 84
rect 52 78 56 82
rect 60 78 64 82
rect 52 76 64 78
rect 67 82 77 84
rect 67 78 71 82
rect 75 78 77 82
rect 67 76 77 78
rect 81 82 91 84
rect 81 78 83 82
rect 87 78 91 82
rect 81 76 91 78
rect 93 82 103 84
rect 93 78 97 82
rect 101 78 103 82
rect 93 76 103 78
rect 428 216 430 220
rect 434 216 438 220
rect 428 214 438 216
rect 441 220 453 222
rect 441 216 445 220
rect 449 216 453 220
rect 441 214 453 216
rect 456 220 466 222
rect 456 216 460 220
rect 464 216 466 220
rect 456 214 466 216
rect 360 172 370 174
rect 360 168 362 172
rect 366 168 370 172
rect 360 166 370 168
rect 373 172 385 174
rect 373 168 377 172
rect 381 168 385 172
rect 373 166 385 168
rect 388 172 398 174
rect 388 168 392 172
rect 396 168 398 172
rect 388 166 398 168
rect 291 82 301 84
rect 291 78 293 82
rect 297 78 301 82
rect 291 76 301 78
rect 304 82 316 84
rect 304 78 308 82
rect 312 78 316 82
rect 304 76 316 78
rect 319 82 329 84
rect 319 78 323 82
rect 327 78 329 82
rect 319 76 329 78
rect 333 82 343 84
rect 333 78 335 82
rect 339 78 343 82
rect 333 76 343 78
rect 345 82 355 84
rect 345 78 349 82
rect 353 78 355 82
rect 345 76 355 78
rect 408 82 418 84
rect 408 78 410 82
rect 414 78 418 82
rect 408 76 418 78
rect 421 76 433 84
rect 436 82 446 84
rect 436 78 440 82
rect 444 78 446 82
rect 436 76 446 78
rect 450 82 460 84
rect 450 78 452 82
rect 456 78 460 82
rect 450 76 460 78
rect 462 82 472 84
rect 462 78 466 82
rect 470 78 472 82
rect 462 76 472 78
rect 877 439 887 441
rect 877 435 879 439
rect 883 435 887 439
rect 877 433 887 435
rect 890 439 902 441
rect 890 435 894 439
rect 898 435 902 439
rect 890 433 902 435
rect 905 439 915 441
rect 905 435 909 439
rect 913 435 915 439
rect 905 433 915 435
rect 810 400 820 402
rect 810 396 812 400
rect 816 396 820 400
rect 810 394 820 396
rect 823 400 835 402
rect 823 396 827 400
rect 831 396 835 400
rect 823 394 835 396
rect 838 400 848 402
rect 945 404 955 406
rect 838 396 842 400
rect 846 396 848 400
rect 838 394 848 396
rect 945 400 947 404
rect 951 400 955 404
rect 945 398 955 400
rect 958 404 970 406
rect 958 400 962 404
rect 966 400 970 404
rect 958 398 970 400
rect 973 404 983 406
rect 973 400 977 404
rect 981 400 983 404
rect 973 398 983 400
rect 877 356 887 358
rect 877 352 879 356
rect 883 352 887 356
rect 877 350 887 352
rect 890 356 902 358
rect 890 352 894 356
rect 898 352 902 356
rect 890 350 902 352
rect 905 356 915 358
rect 905 352 909 356
rect 913 352 915 356
rect 905 350 915 352
rect 648 255 658 257
rect 648 251 650 255
rect 654 251 658 255
rect 648 249 658 251
rect 661 255 673 257
rect 661 251 665 255
rect 669 251 673 255
rect 661 249 673 251
rect 676 255 686 257
rect 676 251 680 255
rect 684 251 686 255
rect 676 249 686 251
rect 883 255 893 257
rect 883 251 885 255
rect 889 251 893 255
rect 883 249 893 251
rect 896 255 908 257
rect 896 251 900 255
rect 904 251 908 255
rect 896 249 908 251
rect 911 255 921 257
rect 911 251 915 255
rect 919 251 921 255
rect 911 249 921 251
rect 581 216 591 218
rect 581 212 583 216
rect 587 212 591 216
rect 581 210 591 212
rect 594 216 606 218
rect 594 212 598 216
rect 602 212 606 216
rect 594 210 606 212
rect 609 216 619 218
rect 716 220 726 222
rect 609 212 613 216
rect 617 212 619 216
rect 609 210 619 212
rect 716 216 718 220
rect 722 216 726 220
rect 716 214 726 216
rect 729 220 741 222
rect 729 216 733 220
rect 737 216 741 220
rect 729 214 741 216
rect 744 220 754 222
rect 744 216 748 220
rect 752 216 754 220
rect 744 214 754 216
rect 816 216 826 218
rect 816 212 818 216
rect 822 212 826 216
rect 816 210 826 212
rect 829 216 841 218
rect 829 212 833 216
rect 837 212 841 216
rect 829 210 841 212
rect 844 216 854 218
rect 951 220 961 222
rect 844 212 848 216
rect 852 212 854 216
rect 844 210 854 212
rect 648 172 658 174
rect 648 168 650 172
rect 654 168 658 172
rect 648 166 658 168
rect 661 172 673 174
rect 661 168 665 172
rect 669 168 673 172
rect 661 166 673 168
rect 676 172 686 174
rect 676 168 680 172
rect 684 168 686 172
rect 676 166 686 168
rect 562 82 572 84
rect 562 78 564 82
rect 568 78 572 82
rect 562 76 572 78
rect 575 82 587 84
rect 575 78 579 82
rect 583 78 587 82
rect 575 76 587 78
rect 590 82 600 84
rect 590 78 594 82
rect 598 78 600 82
rect 590 76 600 78
rect 604 82 614 84
rect 604 78 606 82
rect 610 78 614 82
rect 604 76 614 78
rect 616 82 626 84
rect 616 78 620 82
rect 624 78 626 82
rect 616 76 626 78
rect 951 216 953 220
rect 957 216 961 220
rect 951 214 961 216
rect 964 220 976 222
rect 964 216 968 220
rect 972 216 976 220
rect 964 214 976 216
rect 979 220 989 222
rect 979 216 983 220
rect 987 216 989 220
rect 979 214 989 216
rect 883 172 893 174
rect 883 168 885 172
rect 889 168 893 172
rect 883 166 893 168
rect 896 172 908 174
rect 896 168 900 172
rect 904 168 908 172
rect 896 166 908 168
rect 911 172 921 174
rect 911 168 915 172
rect 919 168 921 172
rect 911 166 921 168
rect 814 82 824 84
rect 814 78 816 82
rect 820 78 824 82
rect 814 76 824 78
rect 827 82 839 84
rect 827 78 831 82
rect 835 78 839 82
rect 827 76 839 78
rect 842 82 852 84
rect 842 78 846 82
rect 850 78 852 82
rect 842 76 852 78
rect 856 82 866 84
rect 856 78 858 82
rect 862 78 866 82
rect 856 76 866 78
rect 868 82 878 84
rect 868 78 872 82
rect 876 78 878 82
rect 868 76 878 78
rect 931 82 941 84
rect 931 78 933 82
rect 937 78 941 82
rect 931 76 941 78
rect 944 76 956 84
rect 959 82 969 84
rect 959 78 963 82
rect 967 78 969 82
rect 959 76 969 78
rect 973 82 983 84
rect 973 78 975 82
rect 979 78 983 82
rect 973 76 983 78
rect 985 82 995 84
rect 985 78 989 82
rect 993 78 995 82
rect 985 76 995 78
rect 1401 439 1411 441
rect 1401 435 1403 439
rect 1407 435 1411 439
rect 1401 433 1411 435
rect 1414 439 1426 441
rect 1414 435 1418 439
rect 1422 435 1426 439
rect 1414 433 1426 435
rect 1429 439 1439 441
rect 1429 435 1433 439
rect 1437 435 1439 439
rect 1429 433 1439 435
rect 1334 400 1344 402
rect 1334 396 1336 400
rect 1340 396 1344 400
rect 1334 394 1344 396
rect 1347 400 1359 402
rect 1347 396 1351 400
rect 1355 396 1359 400
rect 1347 394 1359 396
rect 1362 400 1372 402
rect 1469 404 1479 406
rect 1362 396 1366 400
rect 1370 396 1372 400
rect 1362 394 1372 396
rect 1469 400 1471 404
rect 1475 400 1479 404
rect 1469 398 1479 400
rect 1482 404 1494 406
rect 1482 400 1486 404
rect 1490 400 1494 404
rect 1482 398 1494 400
rect 1497 404 1507 406
rect 1497 400 1501 404
rect 1505 400 1507 404
rect 1497 398 1507 400
rect 1401 356 1411 358
rect 1401 352 1403 356
rect 1407 352 1411 356
rect 1401 350 1411 352
rect 1414 356 1426 358
rect 1414 352 1418 356
rect 1422 352 1426 356
rect 1414 350 1426 352
rect 1429 356 1439 358
rect 1429 352 1433 356
rect 1437 352 1439 356
rect 1429 350 1439 352
rect 1171 255 1181 257
rect 1171 251 1173 255
rect 1177 251 1181 255
rect 1171 249 1181 251
rect 1184 255 1196 257
rect 1184 251 1188 255
rect 1192 251 1196 255
rect 1184 249 1196 251
rect 1199 255 1209 257
rect 1199 251 1203 255
rect 1207 251 1209 255
rect 1199 249 1209 251
rect 1406 255 1416 257
rect 1406 251 1408 255
rect 1412 251 1416 255
rect 1406 249 1416 251
rect 1419 255 1431 257
rect 1419 251 1423 255
rect 1427 251 1431 255
rect 1419 249 1431 251
rect 1434 255 1444 257
rect 1434 251 1438 255
rect 1442 251 1444 255
rect 1434 249 1444 251
rect 1104 216 1114 218
rect 1104 212 1106 216
rect 1110 212 1114 216
rect 1104 210 1114 212
rect 1117 216 1129 218
rect 1117 212 1121 216
rect 1125 212 1129 216
rect 1117 210 1129 212
rect 1132 216 1142 218
rect 1239 220 1249 222
rect 1132 212 1136 216
rect 1140 212 1142 216
rect 1132 210 1142 212
rect 1239 216 1241 220
rect 1245 216 1249 220
rect 1239 214 1249 216
rect 1252 220 1264 222
rect 1252 216 1256 220
rect 1260 216 1264 220
rect 1252 214 1264 216
rect 1267 220 1277 222
rect 1267 216 1271 220
rect 1275 216 1277 220
rect 1267 214 1277 216
rect 1339 216 1349 218
rect 1339 212 1341 216
rect 1345 212 1349 216
rect 1339 210 1349 212
rect 1352 216 1364 218
rect 1352 212 1356 216
rect 1360 212 1364 216
rect 1352 210 1364 212
rect 1367 216 1377 218
rect 1474 220 1484 222
rect 1367 212 1371 216
rect 1375 212 1377 216
rect 1367 210 1377 212
rect 1171 172 1181 174
rect 1171 168 1173 172
rect 1177 168 1181 172
rect 1171 166 1181 168
rect 1184 172 1196 174
rect 1184 168 1188 172
rect 1192 168 1196 172
rect 1184 166 1196 168
rect 1199 172 1209 174
rect 1199 168 1203 172
rect 1207 168 1209 172
rect 1199 166 1209 168
rect 1085 82 1095 84
rect 1085 78 1087 82
rect 1091 78 1095 82
rect 1085 76 1095 78
rect 1098 82 1110 84
rect 1098 78 1102 82
rect 1106 78 1110 82
rect 1098 76 1110 78
rect 1113 82 1123 84
rect 1113 78 1117 82
rect 1121 78 1123 82
rect 1113 76 1123 78
rect 1127 82 1137 84
rect 1127 78 1129 82
rect 1133 78 1137 82
rect 1127 76 1137 78
rect 1139 82 1149 84
rect 1139 78 1143 82
rect 1147 78 1149 82
rect 1139 76 1149 78
rect 1474 216 1476 220
rect 1480 216 1484 220
rect 1474 214 1484 216
rect 1487 220 1499 222
rect 1487 216 1491 220
rect 1495 216 1499 220
rect 1487 214 1499 216
rect 1502 220 1512 222
rect 1502 216 1506 220
rect 1510 216 1512 220
rect 1502 214 1512 216
rect 1406 172 1416 174
rect 1406 168 1408 172
rect 1412 168 1416 172
rect 1406 166 1416 168
rect 1419 172 1431 174
rect 1419 168 1423 172
rect 1427 168 1431 172
rect 1419 166 1431 168
rect 1434 172 1444 174
rect 1434 168 1438 172
rect 1442 168 1444 172
rect 1434 166 1444 168
rect 1337 82 1347 84
rect 1337 78 1339 82
rect 1343 78 1347 82
rect 1337 76 1347 78
rect 1350 82 1362 84
rect 1350 78 1354 82
rect 1358 78 1362 82
rect 1350 76 1362 78
rect 1365 82 1375 84
rect 1365 78 1369 82
rect 1373 78 1375 82
rect 1365 76 1375 78
rect 1379 82 1389 84
rect 1379 78 1381 82
rect 1385 78 1389 82
rect 1379 76 1389 78
rect 1391 82 1401 84
rect 1391 78 1395 82
rect 1399 78 1401 82
rect 1391 76 1401 78
rect 1454 82 1464 84
rect 1454 78 1456 82
rect 1460 78 1464 82
rect 1454 76 1464 78
rect 1467 76 1479 84
rect 1482 82 1492 84
rect 1482 78 1486 82
rect 1490 78 1492 82
rect 1482 76 1492 78
rect 1496 82 1506 84
rect 1496 78 1498 82
rect 1502 78 1506 82
rect 1496 76 1506 78
rect 1508 82 1518 84
rect 1508 78 1512 82
rect 1516 78 1518 82
rect 1508 76 1518 78
rect 1694 255 1704 257
rect 1694 251 1696 255
rect 1700 251 1704 255
rect 1694 249 1704 251
rect 1707 255 1719 257
rect 1707 251 1711 255
rect 1715 251 1719 255
rect 1707 249 1719 251
rect 1722 255 1732 257
rect 1722 251 1726 255
rect 1730 251 1732 255
rect 1722 249 1732 251
rect 1929 255 1939 257
rect 1929 251 1931 255
rect 1935 251 1939 255
rect 1929 249 1939 251
rect 1942 255 1954 257
rect 1942 251 1946 255
rect 1950 251 1954 255
rect 1942 249 1954 251
rect 1957 255 1967 257
rect 1957 251 1961 255
rect 1965 251 1967 255
rect 1957 249 1967 251
rect 1627 216 1637 218
rect 1627 212 1629 216
rect 1633 212 1637 216
rect 1627 210 1637 212
rect 1640 216 1652 218
rect 1640 212 1644 216
rect 1648 212 1652 216
rect 1640 210 1652 212
rect 1655 216 1665 218
rect 1762 220 1772 222
rect 1655 212 1659 216
rect 1663 212 1665 216
rect 1655 210 1665 212
rect 1762 216 1764 220
rect 1768 216 1772 220
rect 1762 214 1772 216
rect 1775 220 1787 222
rect 1775 216 1779 220
rect 1783 216 1787 220
rect 1775 214 1787 216
rect 1790 220 1800 222
rect 1790 216 1794 220
rect 1798 216 1800 220
rect 1790 214 1800 216
rect 1862 216 1872 218
rect 1862 212 1864 216
rect 1868 212 1872 216
rect 1862 210 1872 212
rect 1875 216 1887 218
rect 1875 212 1879 216
rect 1883 212 1887 216
rect 1875 210 1887 212
rect 1890 216 1900 218
rect 1997 220 2007 222
rect 1890 212 1894 216
rect 1898 212 1900 216
rect 1890 210 1900 212
rect 1694 172 1704 174
rect 1694 168 1696 172
rect 1700 168 1704 172
rect 1694 166 1704 168
rect 1707 172 1719 174
rect 1707 168 1711 172
rect 1715 168 1719 172
rect 1707 166 1719 168
rect 1722 172 1732 174
rect 1722 168 1726 172
rect 1730 168 1732 172
rect 1722 166 1732 168
rect 1608 82 1618 84
rect 1608 78 1610 82
rect 1614 78 1618 82
rect 1608 76 1618 78
rect 1621 82 1633 84
rect 1621 78 1625 82
rect 1629 78 1633 82
rect 1621 76 1633 78
rect 1636 82 1646 84
rect 1636 78 1640 82
rect 1644 78 1646 82
rect 1636 76 1646 78
rect 1650 82 1660 84
rect 1650 78 1652 82
rect 1656 78 1660 82
rect 1650 76 1660 78
rect 1662 82 1672 84
rect 1662 78 1666 82
rect 1670 78 1672 82
rect 1662 76 1672 78
rect 1997 216 1999 220
rect 2003 216 2007 220
rect 1997 214 2007 216
rect 2010 220 2022 222
rect 2010 216 2014 220
rect 2018 216 2022 220
rect 2010 214 2022 216
rect 2025 220 2035 222
rect 2025 216 2029 220
rect 2033 216 2035 220
rect 2025 214 2035 216
rect 1929 172 1939 174
rect 1929 168 1931 172
rect 1935 168 1939 172
rect 1929 166 1939 168
rect 1942 172 1954 174
rect 1942 168 1946 172
rect 1950 168 1954 172
rect 1942 166 1954 168
rect 1957 172 1967 174
rect 1957 168 1961 172
rect 1965 168 1967 172
rect 1957 166 1967 168
rect 1860 82 1870 84
rect 1860 78 1862 82
rect 1866 78 1870 82
rect 1860 76 1870 78
rect 1873 82 1885 84
rect 1873 78 1877 82
rect 1881 78 1885 82
rect 1873 76 1885 78
rect 1888 82 1898 84
rect 1888 78 1892 82
rect 1896 78 1898 82
rect 1888 76 1898 78
rect 1902 82 1912 84
rect 1902 78 1904 82
rect 1908 78 1912 82
rect 1902 76 1912 78
rect 1914 82 1924 84
rect 1914 78 1918 82
rect 1922 78 1924 82
rect 1914 76 1924 78
rect 1977 82 1987 84
rect 1977 78 1979 82
rect 1983 78 1987 82
rect 1977 76 1987 78
rect 1990 76 2002 84
rect 2005 82 2015 84
rect 2005 78 2009 82
rect 2013 78 2015 82
rect 2005 76 2015 78
rect 2019 82 2029 84
rect 2019 78 2021 82
rect 2025 78 2029 82
rect 2019 76 2029 78
rect 2031 82 2041 84
rect 2031 78 2035 82
rect 2039 78 2041 82
rect 2031 76 2041 78
<< metal1 >>
rect -232 451 -135 453
rect -232 449 -172 451
rect -168 449 -135 451
rect -131 449 -116 453
rect -112 451 378 453
rect -112 449 341 451
rect -140 439 -136 449
rect -110 439 -106 449
rect -125 426 -121 435
rect -125 422 -106 426
rect -219 418 -144 422
rect -110 418 -106 422
rect -55 418 -51 449
rect 345 449 378 451
rect 382 449 397 453
rect 401 451 884 453
rect 401 449 847 451
rect 373 439 377 449
rect 403 439 407 449
rect 388 426 392 435
rect 388 422 407 426
rect 294 418 369 422
rect 403 418 407 422
rect 458 418 462 449
rect 851 449 884 451
rect 888 449 903 453
rect 907 451 1408 453
rect 907 449 1371 451
rect 879 439 883 449
rect 909 439 913 449
rect 894 426 898 435
rect 894 422 913 426
rect 800 418 875 422
rect 909 418 913 422
rect 964 418 968 449
rect 1375 449 1408 451
rect 1412 449 1427 453
rect 1431 449 2079 453
rect 1403 439 1407 449
rect 1433 439 1437 449
rect 1418 426 1422 435
rect 1418 422 1437 426
rect 1324 418 1399 422
rect 1433 418 1437 422
rect 1488 418 1492 449
rect -219 379 -214 418
rect -148 414 -122 418
rect -110 414 -90 418
rect -74 414 -67 418
rect -63 414 -48 418
rect -44 414 -34 418
rect -211 410 -202 414
rect -198 410 -183 414
rect -179 410 -174 414
rect -207 400 -203 410
rect -177 400 -173 410
rect -157 406 -137 410
rect -192 387 -188 396
rect -192 383 -173 387
rect -177 379 -173 383
rect -157 379 -153 406
rect -110 399 -106 414
rect -140 387 -136 395
rect -142 383 -135 387
rect -131 383 -114 387
rect -110 383 -106 387
rect -94 383 -90 414
rect -72 404 -68 414
rect -42 404 -38 414
rect -57 391 -53 400
rect -57 387 -38 391
rect -42 383 -38 387
rect -94 379 -54 383
rect -42 381 13 383
rect -42 379 9 381
rect -228 375 -189 379
rect -177 375 -153 379
rect -243 367 -204 371
rect -243 287 -239 367
rect -217 340 -212 367
rect -177 360 -173 375
rect -207 348 -203 356
rect -209 344 -202 348
rect -198 344 -181 348
rect -177 344 -172 348
rect -217 336 -162 340
rect -167 327 -162 336
rect -157 335 -153 375
rect -94 371 -69 375
rect -141 366 -135 370
rect -131 366 -116 370
rect -112 366 -104 370
rect -140 356 -136 366
rect -110 356 -106 366
rect -125 343 -121 352
rect -125 339 -106 343
rect -110 335 -106 339
rect -94 335 -90 371
rect -42 364 -38 379
rect 294 379 299 418
rect 365 414 391 418
rect 403 414 423 418
rect 439 414 446 418
rect 450 414 465 418
rect 469 414 479 418
rect 302 410 311 414
rect 315 410 330 414
rect 334 410 339 414
rect 306 400 310 410
rect 336 400 340 410
rect 356 406 376 410
rect 321 387 325 396
rect 321 383 340 387
rect 336 379 340 383
rect 356 379 360 406
rect 403 399 407 414
rect 373 387 377 395
rect 371 383 378 387
rect 382 383 399 387
rect 403 383 407 387
rect 419 383 423 414
rect 441 404 445 414
rect 471 404 475 414
rect 456 391 460 400
rect 456 387 475 391
rect 471 383 475 387
rect 419 379 459 383
rect 471 381 536 383
rect 471 379 532 381
rect 285 375 324 379
rect 336 375 360 379
rect 285 367 309 371
rect -72 352 -68 360
rect -72 348 -67 352
rect -63 348 -46 352
rect -42 348 -38 352
rect 296 340 301 367
rect 336 360 340 375
rect 306 348 310 356
rect 304 344 311 348
rect 315 344 332 348
rect 336 344 341 348
rect 296 336 351 340
rect -157 331 -122 335
rect -110 331 -90 335
rect -167 323 -137 327
rect -110 316 -106 331
rect 346 327 351 336
rect 356 335 360 375
rect 419 371 444 375
rect 372 366 378 370
rect 382 366 397 370
rect 401 366 409 370
rect 373 356 377 366
rect 403 356 407 366
rect 388 343 392 352
rect 388 339 407 343
rect 403 335 407 339
rect 419 335 423 371
rect 471 364 475 379
rect 800 379 805 418
rect 871 414 897 418
rect 909 414 929 418
rect 945 414 952 418
rect 956 414 971 418
rect 975 414 985 418
rect 808 410 817 414
rect 821 410 836 414
rect 840 410 845 414
rect 812 400 816 410
rect 842 400 846 410
rect 862 406 882 410
rect 827 387 831 396
rect 827 383 846 387
rect 842 379 846 383
rect 862 379 866 406
rect 909 399 913 414
rect 879 387 883 395
rect 877 383 884 387
rect 888 383 905 387
rect 909 383 913 387
rect 925 383 929 414
rect 947 404 951 414
rect 977 404 981 414
rect 962 391 966 400
rect 962 387 981 391
rect 977 383 981 387
rect 925 379 965 383
rect 977 381 1059 383
rect 977 379 1055 381
rect 791 375 830 379
rect 842 375 866 379
rect 791 367 815 371
rect 441 352 445 360
rect 441 348 446 352
rect 450 348 467 352
rect 471 348 475 352
rect 802 340 807 367
rect 842 360 846 375
rect 812 348 816 356
rect 810 344 817 348
rect 821 344 838 348
rect 842 344 847 348
rect 802 336 857 340
rect 356 331 391 335
rect 403 331 423 335
rect 346 323 376 327
rect 403 316 407 331
rect 852 327 857 336
rect 862 335 866 375
rect 925 371 950 375
rect 878 366 884 370
rect 888 366 903 370
rect 907 366 915 370
rect 879 356 883 366
rect 909 356 913 366
rect 894 343 898 352
rect 894 339 913 343
rect 909 335 913 339
rect 925 335 929 371
rect 977 364 981 379
rect 1324 379 1329 418
rect 1395 414 1421 418
rect 1433 414 1453 418
rect 1469 414 1476 418
rect 1480 414 1495 418
rect 1499 414 1509 418
rect 1332 410 1341 414
rect 1345 410 1360 414
rect 1364 410 1369 414
rect 1336 400 1340 410
rect 1366 400 1370 410
rect 1386 406 1406 410
rect 1351 387 1355 396
rect 1351 383 1370 387
rect 1366 379 1370 383
rect 1386 379 1390 406
rect 1433 399 1437 414
rect 1403 387 1407 395
rect 1401 383 1408 387
rect 1412 383 1429 387
rect 1433 383 1437 387
rect 1449 383 1453 414
rect 1471 404 1475 414
rect 1501 404 1505 414
rect 1486 391 1490 400
rect 1486 387 1505 391
rect 1501 383 1505 387
rect 1449 379 1489 383
rect 1501 381 1582 383
rect 1501 379 1578 381
rect 1315 375 1354 379
rect 1366 375 1390 379
rect 1315 367 1339 371
rect 947 352 951 360
rect 947 348 952 352
rect 956 348 973 352
rect 977 348 981 352
rect 1326 340 1331 367
rect 1366 360 1370 375
rect 1336 348 1340 356
rect 1334 344 1341 348
rect 1345 344 1362 348
rect 1366 344 1371 348
rect 1326 336 1381 340
rect 862 331 897 335
rect 909 331 929 335
rect 852 323 882 327
rect 909 316 913 331
rect 1376 327 1381 336
rect 1386 335 1390 375
rect 1449 371 1474 375
rect 1402 366 1408 370
rect 1412 366 1427 370
rect 1431 366 1439 370
rect 1403 356 1407 366
rect 1433 356 1437 366
rect 1418 343 1422 352
rect 1418 339 1437 343
rect 1433 335 1437 339
rect 1449 335 1453 371
rect 1501 364 1505 379
rect 1471 352 1475 360
rect 1471 348 1476 352
rect 1480 348 1497 352
rect 1501 348 1505 352
rect 1386 331 1421 335
rect 1433 331 1453 335
rect 1376 323 1406 327
rect 1433 316 1437 331
rect -232 302 -162 304
rect -140 304 -136 312
rect -158 302 -135 304
rect -232 300 -135 302
rect -131 300 -114 304
rect -110 302 -102 304
rect -98 302 -78 304
rect -74 302 351 304
rect 373 304 377 312
rect 355 302 378 304
rect -110 300 -37 302
rect -33 300 378 302
rect 382 300 399 304
rect 403 302 411 304
rect 415 302 435 304
rect 439 302 857 304
rect 879 304 883 312
rect 861 302 884 304
rect 403 300 884 302
rect 888 300 905 304
rect 909 302 917 304
rect 921 302 941 304
rect 945 302 1381 304
rect 1403 304 1407 312
rect 1385 302 1408 304
rect 909 300 1408 302
rect 1412 300 1429 304
rect 1433 302 1441 304
rect 1445 302 1465 304
rect 1469 302 1655 304
rect 1433 300 1655 302
rect -244 285 279 287
rect 283 285 785 287
rect 789 285 1309 287
rect 1313 285 1655 287
rect -244 283 1655 285
rect -165 108 -161 283
rect 2075 269 2079 449
rect -13 267 132 269
rect -13 265 95 267
rect 99 265 132 267
rect 136 265 151 269
rect 155 267 367 269
rect 155 265 330 267
rect 127 255 131 265
rect 157 255 161 265
rect 142 242 146 251
rect 142 238 161 242
rect 48 234 123 238
rect 157 234 161 238
rect 212 234 216 265
rect 334 265 367 267
rect 371 265 386 269
rect 390 267 655 269
rect 390 265 486 267
rect 362 255 366 265
rect 392 255 396 265
rect 377 242 381 251
rect 377 238 396 242
rect 283 234 358 238
rect 392 234 396 238
rect 447 234 451 265
rect 490 265 618 267
rect 622 265 655 267
rect 659 265 674 269
rect 678 267 890 269
rect 678 265 853 267
rect 650 255 654 265
rect 680 255 684 265
rect 665 242 669 251
rect 665 238 684 242
rect 571 234 646 238
rect 680 234 684 238
rect 735 234 739 265
rect 857 265 890 267
rect 894 265 909 269
rect 913 267 1178 269
rect 913 265 1009 267
rect 885 255 889 265
rect 915 255 919 265
rect 900 242 904 251
rect 900 238 919 242
rect 806 234 881 238
rect 915 234 919 238
rect 970 234 974 265
rect 1013 265 1141 267
rect 1145 265 1178 267
rect 1182 265 1197 269
rect 1201 267 1413 269
rect 1201 265 1376 267
rect 1173 255 1177 265
rect 1203 255 1207 265
rect 1188 242 1192 251
rect 1188 238 1207 242
rect 1094 234 1169 238
rect 1203 234 1207 238
rect 1258 234 1262 265
rect 1380 265 1413 267
rect 1417 265 1432 269
rect 1436 267 1701 269
rect 1436 265 1532 267
rect 1408 255 1412 265
rect 1438 255 1442 265
rect 1423 242 1427 251
rect 1423 238 1442 242
rect 1329 234 1404 238
rect 1438 234 1442 238
rect 1493 234 1497 265
rect 1536 265 1664 267
rect 1668 265 1701 267
rect 1705 265 1720 269
rect 1724 267 1936 269
rect 1724 265 1899 267
rect 1696 255 1700 265
rect 1726 255 1730 265
rect 1711 242 1715 251
rect 1711 238 1730 242
rect 1617 234 1692 238
rect 1726 234 1730 238
rect 1781 234 1785 265
rect 1903 265 1936 267
rect 1940 265 1955 269
rect 1959 267 2079 269
rect 1959 265 2055 267
rect 1931 255 1935 265
rect 1961 255 1965 265
rect 1946 242 1950 251
rect 1946 238 1965 242
rect 1852 234 1927 238
rect 1961 234 1965 238
rect 2016 234 2020 265
rect 2059 265 2079 267
rect 13 193 35 195
rect 48 195 53 234
rect 119 230 145 234
rect 157 230 177 234
rect 193 230 200 234
rect 204 230 219 234
rect 223 230 233 234
rect 56 226 65 230
rect 69 226 84 230
rect 88 226 93 230
rect 60 216 64 226
rect 90 216 94 226
rect 110 222 130 226
rect 75 203 79 212
rect 75 199 94 203
rect 90 195 94 199
rect 110 195 114 222
rect 157 215 161 230
rect 127 203 131 211
rect 125 199 132 203
rect 136 199 153 203
rect 157 199 161 203
rect 173 199 177 230
rect 195 220 199 230
rect 225 220 229 230
rect 210 207 214 216
rect 210 203 229 207
rect 225 199 229 203
rect 283 199 288 234
rect 354 230 380 234
rect 392 230 412 234
rect 428 230 435 234
rect 439 230 454 234
rect 458 230 468 234
rect 291 226 300 230
rect 304 226 319 230
rect 323 226 328 230
rect 295 216 299 226
rect 325 216 329 226
rect 345 222 365 226
rect 310 203 314 212
rect 310 199 329 203
rect 173 195 213 199
rect 225 197 288 199
rect 225 195 254 197
rect 39 193 78 195
rect 9 191 78 193
rect 90 191 114 195
rect -1 185 1 187
rect 5 185 63 187
rect -1 183 35 185
rect 39 183 63 185
rect 50 156 55 183
rect 90 176 94 191
rect 60 164 64 172
rect 58 160 65 164
rect 69 160 86 164
rect 90 160 95 164
rect 50 152 105 156
rect 100 143 105 152
rect 110 151 114 191
rect 173 187 198 191
rect 126 182 132 186
rect 136 182 151 186
rect 155 182 163 186
rect 127 172 131 182
rect 157 172 161 182
rect 142 159 146 168
rect 142 155 161 159
rect 157 151 161 155
rect 173 151 177 187
rect 225 180 229 195
rect 258 195 288 197
rect 325 195 329 199
rect 345 195 349 222
rect 392 215 396 230
rect 362 203 366 211
rect 360 199 367 203
rect 371 199 388 203
rect 392 199 396 203
rect 408 199 412 230
rect 430 220 434 230
rect 460 220 464 230
rect 445 207 449 216
rect 445 203 464 207
rect 460 199 464 203
rect 408 195 448 199
rect 460 197 499 199
rect 460 195 495 197
rect 283 191 313 195
rect 325 191 349 195
rect 268 185 298 187
rect 272 183 298 185
rect 195 168 199 176
rect 195 164 200 168
rect 204 164 221 168
rect 225 164 229 168
rect 285 156 290 183
rect 325 176 329 191
rect 295 164 299 172
rect 293 160 300 164
rect 304 160 321 164
rect 325 160 330 164
rect 285 152 340 156
rect 110 147 145 151
rect 157 147 177 151
rect 100 139 130 143
rect 157 132 161 147
rect 335 143 340 152
rect 345 151 349 191
rect 408 187 433 191
rect 361 182 367 186
rect 371 182 386 186
rect 390 182 398 186
rect 362 172 366 182
rect 392 172 396 182
rect 377 159 381 168
rect 377 155 396 159
rect 392 151 396 155
rect 408 151 412 187
rect 460 180 464 195
rect 536 193 558 195
rect 571 195 576 234
rect 642 230 668 234
rect 680 230 700 234
rect 716 230 723 234
rect 727 230 742 234
rect 746 230 756 234
rect 579 226 588 230
rect 592 226 607 230
rect 611 226 616 230
rect 583 216 587 226
rect 613 216 617 226
rect 633 222 653 226
rect 598 203 602 212
rect 598 199 617 203
rect 613 195 617 199
rect 633 195 637 222
rect 680 215 684 230
rect 650 203 654 211
rect 648 199 655 203
rect 659 199 676 203
rect 680 199 684 203
rect 696 199 700 230
rect 718 220 722 230
rect 748 220 752 230
rect 733 207 737 216
rect 733 203 752 207
rect 748 199 752 203
rect 806 199 811 234
rect 877 230 903 234
rect 915 230 935 234
rect 951 230 958 234
rect 962 230 977 234
rect 981 230 991 234
rect 814 226 823 230
rect 827 226 842 230
rect 846 226 851 230
rect 818 216 822 226
rect 848 216 852 226
rect 868 222 888 226
rect 833 203 837 212
rect 833 199 852 203
rect 696 195 736 199
rect 748 197 811 199
rect 748 195 777 197
rect 562 193 601 195
rect 532 191 601 193
rect 613 191 637 195
rect 522 185 524 187
rect 528 185 586 187
rect 522 183 558 185
rect 562 183 586 185
rect 430 168 434 176
rect 430 164 435 168
rect 439 164 456 168
rect 460 164 464 168
rect 573 156 578 183
rect 613 176 617 191
rect 583 164 587 172
rect 581 160 588 164
rect 592 160 609 164
rect 613 160 618 164
rect 573 152 628 156
rect 345 147 380 151
rect 392 147 412 151
rect 335 139 365 143
rect 392 132 396 147
rect 623 143 628 152
rect 633 151 637 191
rect 696 187 721 191
rect 649 182 655 186
rect 659 182 674 186
rect 678 182 686 186
rect 650 172 654 182
rect 680 172 684 182
rect 665 159 669 168
rect 665 155 684 159
rect 680 151 684 155
rect 696 151 700 187
rect 748 180 752 195
rect 781 195 811 197
rect 848 195 852 199
rect 868 195 872 222
rect 915 215 919 230
rect 885 203 889 211
rect 883 199 890 203
rect 894 199 911 203
rect 915 199 919 203
rect 931 199 935 230
rect 953 220 957 230
rect 983 220 987 230
rect 968 207 972 216
rect 968 203 987 207
rect 983 199 987 203
rect 931 195 971 199
rect 983 197 1022 199
rect 983 195 1018 197
rect 806 191 836 195
rect 848 191 872 195
rect 791 185 821 187
rect 795 183 821 185
rect 718 168 722 176
rect 718 164 723 168
rect 727 164 744 168
rect 748 164 752 168
rect 808 156 813 183
rect 848 176 852 191
rect 818 164 822 172
rect 816 160 823 164
rect 827 160 844 164
rect 848 160 853 164
rect 808 152 863 156
rect 633 147 668 151
rect 680 147 700 151
rect 623 139 653 143
rect 680 132 684 147
rect 858 143 863 152
rect 868 151 872 191
rect 931 187 956 191
rect 884 182 890 186
rect 894 182 909 186
rect 913 182 921 186
rect 885 172 889 182
rect 915 172 919 182
rect 900 159 904 168
rect 900 155 919 159
rect 915 151 919 155
rect 931 151 935 187
rect 983 180 987 195
rect 1059 193 1081 195
rect 1094 195 1099 234
rect 1165 230 1191 234
rect 1203 230 1223 234
rect 1239 230 1246 234
rect 1250 230 1265 234
rect 1269 230 1279 234
rect 1102 226 1111 230
rect 1115 226 1130 230
rect 1134 226 1139 230
rect 1106 216 1110 226
rect 1136 216 1140 226
rect 1156 222 1176 226
rect 1121 203 1125 212
rect 1121 199 1140 203
rect 1136 195 1140 199
rect 1156 195 1160 222
rect 1203 215 1207 230
rect 1173 203 1177 211
rect 1171 199 1178 203
rect 1182 199 1199 203
rect 1203 199 1207 203
rect 1219 199 1223 230
rect 1241 220 1245 230
rect 1271 220 1275 230
rect 1256 207 1260 216
rect 1256 203 1275 207
rect 1271 199 1275 203
rect 1329 199 1334 234
rect 1400 230 1426 234
rect 1438 230 1458 234
rect 1474 230 1481 234
rect 1485 230 1500 234
rect 1504 230 1514 234
rect 1337 226 1346 230
rect 1350 226 1365 230
rect 1369 226 1374 230
rect 1341 216 1345 226
rect 1371 216 1375 226
rect 1391 222 1411 226
rect 1356 203 1360 212
rect 1356 199 1375 203
rect 1219 195 1259 199
rect 1271 197 1334 199
rect 1271 195 1300 197
rect 1085 193 1124 195
rect 1055 191 1124 193
rect 1136 191 1160 195
rect 1045 185 1047 187
rect 1051 185 1109 187
rect 1045 183 1081 185
rect 1085 183 1109 185
rect 953 168 957 176
rect 953 164 958 168
rect 962 164 979 168
rect 983 164 987 168
rect 1096 156 1101 183
rect 1136 176 1140 191
rect 1106 164 1110 172
rect 1104 160 1111 164
rect 1115 160 1132 164
rect 1136 160 1141 164
rect 1096 152 1151 156
rect 868 147 903 151
rect 915 147 935 151
rect 858 139 888 143
rect 915 132 919 147
rect 1146 143 1151 152
rect 1156 151 1160 191
rect 1219 187 1244 191
rect 1172 182 1178 186
rect 1182 182 1197 186
rect 1201 182 1209 186
rect 1173 172 1177 182
rect 1203 172 1207 182
rect 1188 159 1192 168
rect 1188 155 1207 159
rect 1203 151 1207 155
rect 1219 151 1223 187
rect 1271 180 1275 195
rect 1304 195 1334 197
rect 1371 195 1375 199
rect 1391 195 1395 222
rect 1438 215 1442 230
rect 1408 203 1412 211
rect 1406 199 1413 203
rect 1417 199 1434 203
rect 1438 199 1442 203
rect 1454 199 1458 230
rect 1476 220 1480 230
rect 1506 220 1510 230
rect 1491 207 1495 216
rect 1491 203 1510 207
rect 1506 199 1510 203
rect 1454 195 1494 199
rect 1506 197 1545 199
rect 1506 195 1541 197
rect 1329 191 1359 195
rect 1371 191 1395 195
rect 1314 185 1344 187
rect 1318 183 1344 185
rect 1241 168 1245 176
rect 1241 164 1246 168
rect 1250 164 1267 168
rect 1271 164 1275 168
rect 1331 156 1336 183
rect 1371 176 1375 191
rect 1341 164 1345 172
rect 1339 160 1346 164
rect 1350 160 1367 164
rect 1371 160 1376 164
rect 1331 152 1386 156
rect 1156 147 1191 151
rect 1203 147 1223 151
rect 1146 139 1176 143
rect 1203 132 1207 147
rect 1381 143 1386 152
rect 1391 151 1395 191
rect 1454 187 1479 191
rect 1407 182 1413 186
rect 1417 182 1432 186
rect 1436 182 1444 186
rect 1408 172 1412 182
rect 1438 172 1442 182
rect 1423 159 1427 168
rect 1423 155 1442 159
rect 1438 151 1442 155
rect 1454 151 1458 187
rect 1506 180 1510 195
rect 1582 193 1604 195
rect 1617 195 1622 234
rect 1688 230 1714 234
rect 1726 230 1746 234
rect 1762 230 1769 234
rect 1773 230 1788 234
rect 1792 230 1802 234
rect 1625 226 1634 230
rect 1638 226 1653 230
rect 1657 226 1662 230
rect 1629 216 1633 226
rect 1659 216 1663 226
rect 1679 222 1699 226
rect 1644 203 1648 212
rect 1644 199 1663 203
rect 1659 195 1663 199
rect 1679 195 1683 222
rect 1726 215 1730 230
rect 1696 203 1700 211
rect 1694 199 1701 203
rect 1705 199 1722 203
rect 1726 199 1730 203
rect 1742 199 1746 230
rect 1764 220 1768 230
rect 1794 220 1798 230
rect 1779 207 1783 216
rect 1779 203 1798 207
rect 1794 199 1798 203
rect 1852 199 1857 234
rect 1923 230 1949 234
rect 1961 230 1981 234
rect 1997 230 2004 234
rect 2008 230 2023 234
rect 2027 230 2037 234
rect 1860 226 1869 230
rect 1873 226 1888 230
rect 1892 226 1897 230
rect 1864 216 1868 226
rect 1894 216 1898 226
rect 1914 222 1934 226
rect 1879 203 1883 212
rect 1879 199 1898 203
rect 1742 195 1782 199
rect 1794 197 1857 199
rect 1794 195 1823 197
rect 1608 193 1647 195
rect 1578 191 1647 193
rect 1659 191 1683 195
rect 1568 185 1570 187
rect 1574 185 1632 187
rect 1568 183 1604 185
rect 1608 183 1632 185
rect 1476 168 1480 176
rect 1476 164 1481 168
rect 1485 164 1502 168
rect 1506 164 1510 168
rect 1619 156 1624 183
rect 1659 176 1663 191
rect 1629 164 1633 172
rect 1627 160 1634 164
rect 1638 160 1655 164
rect 1659 160 1664 164
rect 1619 152 1674 156
rect 1391 147 1426 151
rect 1438 147 1458 151
rect 1381 139 1411 143
rect 1438 132 1442 147
rect 1669 143 1674 152
rect 1679 151 1683 191
rect 1742 187 1767 191
rect 1695 182 1701 186
rect 1705 182 1720 186
rect 1724 182 1732 186
rect 1696 172 1700 182
rect 1726 172 1730 182
rect 1711 159 1715 168
rect 1711 155 1730 159
rect 1726 151 1730 155
rect 1742 151 1746 187
rect 1794 180 1798 195
rect 1827 195 1857 197
rect 1894 195 1898 199
rect 1914 195 1918 222
rect 1961 215 1965 230
rect 1931 203 1935 211
rect 1929 199 1936 203
rect 1940 199 1957 203
rect 1961 199 1965 203
rect 1977 199 1981 230
rect 1999 220 2003 230
rect 2029 220 2033 230
rect 2014 207 2018 216
rect 2014 203 2033 207
rect 2029 199 2033 203
rect 1977 195 2017 199
rect 2029 197 2068 199
rect 2029 195 2064 197
rect 1852 191 1882 195
rect 1894 191 1918 195
rect 1837 185 1867 187
rect 1841 183 1867 185
rect 1764 168 1768 176
rect 1764 164 1769 168
rect 1773 164 1790 168
rect 1794 164 1798 168
rect 1854 156 1859 183
rect 1894 176 1898 191
rect 1864 164 1868 172
rect 1862 160 1869 164
rect 1873 160 1890 164
rect 1894 160 1899 164
rect 1854 152 1909 156
rect 1679 147 1714 151
rect 1726 147 1746 151
rect 1669 139 1699 143
rect 1726 132 1730 147
rect 1904 143 1909 152
rect 1914 151 1918 191
rect 1977 187 2002 191
rect 1930 182 1936 186
rect 1940 182 1955 186
rect 1959 182 1967 186
rect 1931 172 1935 182
rect 1961 172 1965 182
rect 1946 159 1950 168
rect 1946 155 1965 159
rect 1961 151 1965 155
rect 1977 151 1981 187
rect 2029 180 2033 195
rect 1999 168 2003 176
rect 1999 164 2004 168
rect 2008 164 2025 168
rect 2029 164 2033 168
rect 1914 147 1949 151
rect 1961 147 1981 151
rect 1904 139 1934 143
rect 1961 132 1965 147
rect 94 118 105 120
rect 127 120 131 128
rect 109 118 132 120
rect 94 116 132 118
rect 136 116 153 120
rect 157 118 165 120
rect 169 118 189 120
rect 193 118 340 120
rect 362 120 366 128
rect 344 118 367 120
rect 157 116 367 118
rect 371 116 388 120
rect 392 118 400 120
rect 404 118 424 120
rect 428 118 492 120
rect 392 116 478 118
rect 482 116 492 118
rect 617 118 628 120
rect 650 120 654 128
rect 632 118 655 120
rect 617 116 655 118
rect 659 116 676 120
rect 680 118 688 120
rect 692 118 712 120
rect 716 118 863 120
rect 885 120 889 128
rect 867 118 890 120
rect 680 116 890 118
rect 894 116 911 120
rect 915 118 923 120
rect 927 118 947 120
rect 951 118 1015 120
rect 915 116 1001 118
rect 1005 116 1015 118
rect 1140 118 1151 120
rect 1173 120 1177 128
rect 1155 118 1178 120
rect 1140 116 1178 118
rect 1182 116 1199 120
rect 1203 118 1211 120
rect 1215 118 1235 120
rect 1239 118 1386 120
rect 1408 120 1412 128
rect 1390 118 1413 120
rect 1203 116 1413 118
rect 1417 116 1434 120
rect 1438 118 1446 120
rect 1450 118 1470 120
rect 1474 118 1538 120
rect 1438 116 1524 118
rect 1528 116 1538 118
rect 1663 118 1674 120
rect 1696 120 1700 128
rect 1678 118 1701 120
rect 1663 116 1701 118
rect 1705 116 1722 120
rect 1726 118 1734 120
rect 1738 118 1758 120
rect 1762 118 1909 120
rect 1931 120 1935 128
rect 1913 118 1936 120
rect 1726 116 1936 118
rect 1940 116 1957 120
rect 1961 118 1969 120
rect 1973 118 1993 120
rect 1997 118 2061 120
rect 1961 116 2047 118
rect 2051 116 2061 118
rect -165 106 268 108
rect -165 104 242 106
rect 246 104 272 106
rect 521 106 791 108
rect 521 104 765 106
rect 38 92 46 96
rect 50 92 65 96
rect 69 92 83 96
rect 87 92 97 96
rect 101 92 298 96
rect 302 92 317 96
rect 321 92 335 96
rect 339 92 349 96
rect 353 92 415 96
rect 419 92 434 96
rect 438 92 452 96
rect 456 92 466 96
rect 470 94 486 96
rect 490 94 492 96
rect 470 92 492 94
rect 41 82 45 92
rect 71 82 75 92
rect 83 82 87 92
rect 293 82 297 92
rect 323 82 327 92
rect 335 82 339 92
rect 410 82 414 92
rect 452 82 456 92
rect 56 69 60 78
rect 56 65 75 69
rect 71 61 75 65
rect 97 63 101 78
rect 308 69 312 78
rect 349 69 353 78
rect 260 65 300 69
rect 308 65 327 69
rect 71 57 87 61
rect 97 59 103 63
rect 296 61 300 65
rect 323 61 327 65
rect 349 65 429 69
rect 71 42 75 57
rect 97 42 101 59
rect 296 57 311 61
rect 323 57 339 61
rect 248 49 296 53
rect 323 42 327 57
rect 349 42 353 65
rect 440 61 444 78
rect 466 63 470 78
rect 521 63 525 104
rect 769 104 795 106
rect 1044 106 1314 108
rect 1044 104 1288 106
rect 561 92 569 96
rect 573 92 588 96
rect 592 92 606 96
rect 610 92 620 96
rect 624 92 821 96
rect 825 92 840 96
rect 844 92 858 96
rect 862 92 872 96
rect 876 92 938 96
rect 942 92 957 96
rect 961 92 975 96
rect 979 92 989 96
rect 993 94 1009 96
rect 1013 94 1015 96
rect 993 92 1015 94
rect 564 82 568 92
rect 594 82 598 92
rect 606 82 610 92
rect 816 82 820 92
rect 846 82 850 92
rect 858 82 862 92
rect 933 82 937 92
rect 975 82 979 92
rect 579 69 583 78
rect 579 65 598 69
rect 424 57 456 61
rect 466 59 525 63
rect 594 61 598 65
rect 620 63 624 78
rect 831 69 835 78
rect 872 69 876 78
rect 783 65 823 69
rect 831 65 850 69
rect 406 49 413 53
rect 424 42 428 57
rect 466 42 470 59
rect 594 57 610 61
rect 620 59 626 63
rect 819 61 823 65
rect 846 61 850 65
rect 872 65 952 69
rect 594 42 598 57
rect 620 42 624 59
rect 819 57 834 61
rect 846 57 862 61
rect 771 49 819 53
rect 846 42 850 57
rect 872 42 876 65
rect 963 61 967 78
rect 989 63 993 78
rect 1044 63 1048 104
rect 1292 104 1318 106
rect 1567 106 1837 108
rect 1567 104 1811 106
rect 1084 92 1092 96
rect 1096 92 1111 96
rect 1115 92 1129 96
rect 1133 92 1143 96
rect 1147 92 1344 96
rect 1348 92 1363 96
rect 1367 92 1381 96
rect 1385 92 1395 96
rect 1399 92 1461 96
rect 1465 92 1480 96
rect 1484 92 1498 96
rect 1502 92 1512 96
rect 1516 94 1532 96
rect 1536 94 1538 96
rect 1516 92 1538 94
rect 1087 82 1091 92
rect 1117 82 1121 92
rect 1129 82 1133 92
rect 1339 82 1343 92
rect 1369 82 1373 92
rect 1381 82 1385 92
rect 1456 82 1460 92
rect 1498 82 1502 92
rect 1102 69 1106 78
rect 1102 65 1121 69
rect 947 57 979 61
rect 989 59 1048 63
rect 1117 61 1121 65
rect 1143 63 1147 78
rect 1354 69 1358 78
rect 1395 69 1399 78
rect 1306 65 1346 69
rect 1354 65 1373 69
rect 929 49 936 53
rect 947 42 951 57
rect 989 42 993 59
rect 1117 57 1133 61
rect 1143 59 1149 63
rect 1342 61 1346 65
rect 1369 61 1373 65
rect 1395 65 1475 69
rect 1117 42 1121 57
rect 1143 42 1147 59
rect 1342 57 1357 61
rect 1369 57 1385 61
rect 1294 49 1342 53
rect 1369 42 1373 57
rect 1395 42 1399 65
rect 1486 61 1490 78
rect 1512 63 1516 78
rect 1567 63 1571 104
rect 1815 104 1841 106
rect 1607 92 1615 96
rect 1619 92 1634 96
rect 1638 92 1652 96
rect 1656 92 1666 96
rect 1670 92 1867 96
rect 1871 92 1886 96
rect 1890 92 1904 96
rect 1908 92 1918 96
rect 1922 92 1984 96
rect 1988 92 2003 96
rect 2007 92 2021 96
rect 2025 92 2035 96
rect 2039 94 2055 96
rect 2059 94 2061 96
rect 2039 92 2061 94
rect 1610 82 1614 92
rect 1640 82 1644 92
rect 1652 82 1656 92
rect 1862 82 1866 92
rect 1892 82 1896 92
rect 1904 82 1908 92
rect 1979 82 1983 92
rect 2021 82 2025 92
rect 1625 69 1629 78
rect 1625 65 1644 69
rect 1470 57 1502 61
rect 1512 59 1571 63
rect 1640 61 1644 65
rect 1666 63 1670 78
rect 1877 69 1881 78
rect 1918 69 1922 78
rect 1829 65 1869 69
rect 1877 65 1896 69
rect 1452 49 1459 53
rect 1470 42 1474 57
rect 1512 42 1516 59
rect 1640 57 1656 61
rect 1666 59 1672 63
rect 1865 61 1869 65
rect 1892 61 1896 65
rect 1918 65 1998 69
rect 1640 42 1644 57
rect 1666 42 1670 59
rect 1865 57 1880 61
rect 1892 57 1908 61
rect 1817 49 1865 53
rect 1892 42 1896 57
rect 1918 42 1922 65
rect 2009 61 2013 78
rect 2035 63 2039 78
rect 1993 57 2025 61
rect 2035 59 2079 63
rect 1975 49 1982 53
rect 1993 42 1997 57
rect 2035 42 2039 59
rect 41 30 45 38
rect 83 30 87 38
rect 293 30 297 38
rect 335 30 339 38
rect 410 30 414 38
rect 440 30 444 38
rect 452 30 456 38
rect -9 28 46 30
rect -13 26 46 28
rect 50 26 67 30
rect 71 26 83 30
rect 87 26 98 30
rect 102 26 298 30
rect 302 26 319 30
rect 323 26 335 30
rect 339 26 350 30
rect 354 26 415 30
rect 419 26 436 30
rect 440 26 452 30
rect 456 26 467 30
rect 471 28 478 30
rect 564 30 568 38
rect 606 30 610 38
rect 816 30 820 38
rect 858 30 862 38
rect 933 30 937 38
rect 963 30 967 38
rect 975 30 979 38
rect 482 28 569 30
rect 471 26 569 28
rect 573 26 590 30
rect 594 26 606 30
rect 610 26 621 30
rect 625 26 821 30
rect 825 26 842 30
rect 846 26 858 30
rect 862 26 873 30
rect 877 26 938 30
rect 942 26 959 30
rect 963 26 975 30
rect 979 26 990 30
rect 994 28 1001 30
rect 1087 30 1091 38
rect 1129 30 1133 38
rect 1339 30 1343 38
rect 1381 30 1385 38
rect 1456 30 1460 38
rect 1486 30 1490 38
rect 1498 30 1502 38
rect 1005 28 1092 30
rect 994 26 1092 28
rect 1096 26 1113 30
rect 1117 26 1129 30
rect 1133 26 1144 30
rect 1148 26 1344 30
rect 1348 26 1365 30
rect 1369 26 1381 30
rect 1385 26 1396 30
rect 1400 26 1461 30
rect 1465 26 1482 30
rect 1486 26 1498 30
rect 1502 26 1513 30
rect 1517 28 1524 30
rect 1610 30 1614 38
rect 1652 30 1656 38
rect 1862 30 1866 38
rect 1904 30 1908 38
rect 1979 30 1983 38
rect 2009 30 2013 38
rect 2021 30 2025 38
rect 1528 28 1615 30
rect 1517 26 1615 28
rect 1619 26 1636 30
rect 1640 26 1652 30
rect 1656 26 1667 30
rect 1671 26 1867 30
rect 1871 26 1888 30
rect 1892 26 1904 30
rect 1908 26 1919 30
rect 1923 26 1984 30
rect 1988 26 2005 30
rect 2009 26 2021 30
rect 2025 26 2036 30
rect 2040 28 2047 30
rect 2051 28 2079 30
rect 2040 26 2079 28
<< metal2 >>
rect -172 414 -168 447
rect 341 414 345 447
rect 847 414 851 447
rect 1371 414 1375 447
rect -170 410 -160 414
rect 343 410 353 414
rect 849 410 859 414
rect 1373 410 1383 414
rect -164 370 -160 410
rect -164 366 -145 370
rect -168 344 -158 348
rect -162 306 -158 344
rect -102 306 -98 387
rect 349 370 353 410
rect 349 366 368 370
rect -78 348 -76 352
rect -78 306 -74 348
rect 345 344 355 348
rect 351 306 355 344
rect 411 306 415 387
rect 855 370 859 410
rect 855 366 874 370
rect 435 348 437 352
rect 435 306 439 348
rect 851 344 861 348
rect 857 306 861 344
rect 917 306 921 387
rect 1379 370 1383 410
rect 1379 366 1398 370
rect 941 348 943 352
rect 941 306 945 348
rect 1375 344 1385 348
rect 1381 306 1385 344
rect 1441 306 1445 387
rect 1465 348 1467 352
rect 1465 306 1469 348
rect -37 160 -33 298
rect 95 230 99 263
rect 330 230 334 263
rect 97 226 107 230
rect 332 226 342 230
rect 103 186 107 226
rect 103 182 122 186
rect 99 160 109 164
rect -37 156 -9 160
rect -13 32 -9 156
rect 105 122 109 160
rect 165 122 169 203
rect 338 186 342 226
rect 338 182 357 186
rect 189 164 191 168
rect 189 122 193 164
rect 334 160 344 164
rect 340 122 344 160
rect 400 122 404 203
rect 424 164 426 168
rect 424 122 428 164
rect 478 32 482 114
rect 486 98 490 263
rect 618 230 622 263
rect 853 230 857 263
rect 620 226 630 230
rect 855 226 865 230
rect 626 186 630 226
rect 626 182 645 186
rect 622 160 632 164
rect 628 122 632 160
rect 688 122 692 203
rect 861 186 865 226
rect 861 182 880 186
rect 712 164 714 168
rect 712 122 716 164
rect 857 160 867 164
rect 863 122 867 160
rect 923 122 927 203
rect 947 164 949 168
rect 947 122 951 164
rect 1001 32 1005 114
rect 1009 98 1013 263
rect 1141 230 1145 263
rect 1376 230 1380 263
rect 1143 226 1153 230
rect 1378 226 1388 230
rect 1149 186 1153 226
rect 1149 182 1168 186
rect 1145 160 1155 164
rect 1151 122 1155 160
rect 1211 122 1215 203
rect 1384 186 1388 226
rect 1384 182 1403 186
rect 1235 164 1237 168
rect 1235 122 1239 164
rect 1380 160 1390 164
rect 1386 122 1390 160
rect 1446 122 1450 203
rect 1470 164 1472 168
rect 1470 122 1474 164
rect 1524 32 1528 114
rect 1532 98 1536 263
rect 1664 230 1668 263
rect 1899 230 1903 263
rect 1666 226 1676 230
rect 1901 226 1911 230
rect 1672 186 1676 226
rect 1672 182 1691 186
rect 1668 160 1678 164
rect 1674 122 1678 160
rect 1734 122 1738 203
rect 1907 186 1911 226
rect 1907 182 1926 186
rect 1758 164 1760 168
rect 1758 122 1762 164
rect 1903 160 1913 164
rect 1909 122 1913 160
rect 1969 122 1973 203
rect 1993 164 1995 168
rect 1993 122 1997 164
rect 2047 32 2051 114
rect 2055 98 2059 263
<< ntransistor >>
rect -132 393 -129 401
rect -117 393 -114 401
rect -199 354 -196 362
rect -184 354 -181 362
rect -64 358 -61 366
rect -49 358 -46 366
rect -132 310 -129 318
rect -117 310 -114 318
rect 381 393 384 401
rect 396 393 399 401
rect 314 354 317 362
rect 329 354 332 362
rect 449 358 452 366
rect 464 358 467 366
rect 381 310 384 318
rect 396 310 399 318
rect 135 209 138 217
rect 150 209 153 217
rect 68 170 71 178
rect 83 170 86 178
rect 203 174 206 182
rect 218 174 221 182
rect 135 126 138 134
rect 150 126 153 134
rect 49 36 52 44
rect 64 36 67 44
rect 91 36 93 44
rect 370 209 373 217
rect 385 209 388 217
rect 303 170 306 178
rect 318 170 321 178
rect 438 174 441 182
rect 453 174 456 182
rect 370 126 373 134
rect 385 126 388 134
rect 301 36 304 44
rect 316 36 319 44
rect 343 36 345 44
rect 418 36 421 44
rect 433 36 436 44
rect 460 36 462 44
rect 887 393 890 401
rect 902 393 905 401
rect 820 354 823 362
rect 835 354 838 362
rect 955 358 958 366
rect 970 358 973 366
rect 887 310 890 318
rect 902 310 905 318
rect 658 209 661 217
rect 673 209 676 217
rect 591 170 594 178
rect 606 170 609 178
rect 726 174 729 182
rect 741 174 744 182
rect 658 126 661 134
rect 673 126 676 134
rect 572 36 575 44
rect 587 36 590 44
rect 614 36 616 44
rect 893 209 896 217
rect 908 209 911 217
rect 826 170 829 178
rect 841 170 844 178
rect 961 174 964 182
rect 976 174 979 182
rect 893 126 896 134
rect 908 126 911 134
rect 824 36 827 44
rect 839 36 842 44
rect 866 36 868 44
rect 941 36 944 44
rect 956 36 959 44
rect 983 36 985 44
rect 1411 393 1414 401
rect 1426 393 1429 401
rect 1344 354 1347 362
rect 1359 354 1362 362
rect 1479 358 1482 366
rect 1494 358 1497 366
rect 1411 310 1414 318
rect 1426 310 1429 318
rect 1181 209 1184 217
rect 1196 209 1199 217
rect 1114 170 1117 178
rect 1129 170 1132 178
rect 1249 174 1252 182
rect 1264 174 1267 182
rect 1181 126 1184 134
rect 1196 126 1199 134
rect 1095 36 1098 44
rect 1110 36 1113 44
rect 1137 36 1139 44
rect 1416 209 1419 217
rect 1431 209 1434 217
rect 1349 170 1352 178
rect 1364 170 1367 178
rect 1484 174 1487 182
rect 1499 174 1502 182
rect 1416 126 1419 134
rect 1431 126 1434 134
rect 1347 36 1350 44
rect 1362 36 1365 44
rect 1389 36 1391 44
rect 1464 36 1467 44
rect 1479 36 1482 44
rect 1506 36 1508 44
rect 1704 209 1707 217
rect 1719 209 1722 217
rect 1637 170 1640 178
rect 1652 170 1655 178
rect 1772 174 1775 182
rect 1787 174 1790 182
rect 1704 126 1707 134
rect 1719 126 1722 134
rect 1618 36 1621 44
rect 1633 36 1636 44
rect 1660 36 1662 44
rect 1939 209 1942 217
rect 1954 209 1957 217
rect 1872 170 1875 178
rect 1887 170 1890 178
rect 2007 174 2010 182
rect 2022 174 2025 182
rect 1939 126 1942 134
rect 1954 126 1957 134
rect 1870 36 1873 44
rect 1885 36 1888 44
rect 1912 36 1914 44
rect 1987 36 1990 44
rect 2002 36 2005 44
rect 2029 36 2031 44
<< ptransistor >>
rect -132 433 -129 441
rect -117 433 -114 441
rect -199 394 -196 402
rect -184 394 -181 402
rect -64 398 -61 406
rect -49 398 -46 406
rect -132 350 -129 358
rect -117 350 -114 358
rect 381 433 384 441
rect 396 433 399 441
rect 314 394 317 402
rect 329 394 332 402
rect 449 398 452 406
rect 464 398 467 406
rect 381 350 384 358
rect 396 350 399 358
rect 135 249 138 257
rect 150 249 153 257
rect 370 249 373 257
rect 385 249 388 257
rect 68 210 71 218
rect 83 210 86 218
rect 203 214 206 222
rect 218 214 221 222
rect 303 210 306 218
rect 318 210 321 218
rect 135 166 138 174
rect 150 166 153 174
rect 49 76 52 84
rect 64 76 67 84
rect 91 76 93 84
rect 438 214 441 222
rect 453 214 456 222
rect 370 166 373 174
rect 385 166 388 174
rect 301 76 304 84
rect 316 76 319 84
rect 343 76 345 84
rect 418 76 421 84
rect 433 76 436 84
rect 460 76 462 84
rect 887 433 890 441
rect 902 433 905 441
rect 820 394 823 402
rect 835 394 838 402
rect 955 398 958 406
rect 970 398 973 406
rect 887 350 890 358
rect 902 350 905 358
rect 658 249 661 257
rect 673 249 676 257
rect 893 249 896 257
rect 908 249 911 257
rect 591 210 594 218
rect 606 210 609 218
rect 726 214 729 222
rect 741 214 744 222
rect 826 210 829 218
rect 841 210 844 218
rect 658 166 661 174
rect 673 166 676 174
rect 572 76 575 84
rect 587 76 590 84
rect 614 76 616 84
rect 961 214 964 222
rect 976 214 979 222
rect 893 166 896 174
rect 908 166 911 174
rect 824 76 827 84
rect 839 76 842 84
rect 866 76 868 84
rect 941 76 944 84
rect 956 76 959 84
rect 983 76 985 84
rect 1411 433 1414 441
rect 1426 433 1429 441
rect 1344 394 1347 402
rect 1359 394 1362 402
rect 1479 398 1482 406
rect 1494 398 1497 406
rect 1411 350 1414 358
rect 1426 350 1429 358
rect 1181 249 1184 257
rect 1196 249 1199 257
rect 1416 249 1419 257
rect 1431 249 1434 257
rect 1114 210 1117 218
rect 1129 210 1132 218
rect 1249 214 1252 222
rect 1264 214 1267 222
rect 1349 210 1352 218
rect 1364 210 1367 218
rect 1181 166 1184 174
rect 1196 166 1199 174
rect 1095 76 1098 84
rect 1110 76 1113 84
rect 1137 76 1139 84
rect 1484 214 1487 222
rect 1499 214 1502 222
rect 1416 166 1419 174
rect 1431 166 1434 174
rect 1347 76 1350 84
rect 1362 76 1365 84
rect 1389 76 1391 84
rect 1464 76 1467 84
rect 1479 76 1482 84
rect 1506 76 1508 84
rect 1704 249 1707 257
rect 1719 249 1722 257
rect 1939 249 1942 257
rect 1954 249 1957 257
rect 1637 210 1640 218
rect 1652 210 1655 218
rect 1772 214 1775 222
rect 1787 214 1790 222
rect 1872 210 1875 218
rect 1887 210 1890 218
rect 1704 166 1707 174
rect 1719 166 1722 174
rect 1618 76 1621 84
rect 1633 76 1636 84
rect 1660 76 1662 84
rect 2007 214 2010 222
rect 2022 214 2025 222
rect 1939 166 1942 174
rect 1954 166 1957 174
rect 1870 76 1873 84
rect 1885 76 1888 84
rect 1912 76 1914 84
rect 1987 76 1990 84
rect 2002 76 2005 84
rect 2029 76 2031 84
<< polycontact >>
rect -122 414 -118 418
rect -137 406 -133 410
rect -232 375 -228 379
rect -189 375 -185 379
rect -54 379 -50 383
rect -204 367 -200 371
rect -69 371 -65 375
rect -122 331 -118 335
rect -137 323 -133 327
rect 9 377 13 381
rect 391 414 395 418
rect 376 406 380 410
rect 281 375 285 379
rect 324 375 328 379
rect 459 379 463 383
rect 281 367 285 371
rect 309 367 313 371
rect 444 371 448 375
rect 391 331 395 335
rect 376 323 380 327
rect 279 285 283 289
rect 145 230 149 234
rect 130 222 134 226
rect 380 230 384 234
rect 365 222 369 226
rect 9 193 13 197
rect 1 185 5 189
rect 35 193 39 197
rect 78 191 82 195
rect 213 195 217 199
rect 35 181 39 185
rect 63 183 67 187
rect 198 187 202 191
rect 254 193 258 197
rect 145 147 149 151
rect 130 139 134 143
rect 242 102 246 106
rect 87 57 91 61
rect 103 59 107 63
rect 313 191 317 195
rect 448 195 452 199
rect 268 181 272 185
rect 298 183 302 187
rect 433 187 437 191
rect 495 193 499 197
rect 380 147 384 151
rect 365 139 369 143
rect 268 106 272 110
rect 256 65 260 69
rect 311 57 315 61
rect 339 57 343 61
rect 244 49 248 53
rect 296 49 300 53
rect 429 65 433 69
rect 413 49 417 53
rect 456 57 460 61
rect 532 377 536 381
rect 897 414 901 418
rect 882 406 886 410
rect 787 375 791 379
rect 830 375 834 379
rect 965 379 969 383
rect 787 367 791 371
rect 815 367 819 371
rect 950 371 954 375
rect 897 331 901 335
rect 882 323 886 327
rect 785 285 789 289
rect 668 230 672 234
rect 653 222 657 226
rect 903 230 907 234
rect 888 222 892 226
rect 532 193 536 197
rect 524 185 528 189
rect 558 193 562 197
rect 601 191 605 195
rect 736 195 740 199
rect 558 181 562 185
rect 586 183 590 187
rect 721 187 725 191
rect 777 193 781 197
rect 668 147 672 151
rect 653 139 657 143
rect 765 102 769 106
rect 610 57 614 61
rect 626 59 630 63
rect 836 191 840 195
rect 971 195 975 199
rect 791 181 795 185
rect 821 183 825 187
rect 956 187 960 191
rect 1018 193 1022 197
rect 903 147 907 151
rect 888 139 892 143
rect 791 106 795 110
rect 779 65 783 69
rect 834 57 838 61
rect 862 57 866 61
rect 767 49 771 53
rect 819 49 823 53
rect 952 65 956 69
rect 936 49 940 53
rect 979 57 983 61
rect 1055 377 1059 381
rect 1421 414 1425 418
rect 1406 406 1410 410
rect 1311 375 1315 379
rect 1354 375 1358 379
rect 1489 379 1493 383
rect 1311 367 1315 371
rect 1339 367 1343 371
rect 1474 371 1478 375
rect 1421 331 1425 335
rect 1406 323 1410 327
rect 1309 285 1313 289
rect 1191 230 1195 234
rect 1176 222 1180 226
rect 1426 230 1430 234
rect 1411 222 1415 226
rect 1055 193 1059 197
rect 1047 185 1051 189
rect 1081 193 1085 197
rect 1124 191 1128 195
rect 1259 195 1263 199
rect 1081 181 1085 185
rect 1109 183 1113 187
rect 1244 187 1248 191
rect 1300 193 1304 197
rect 1191 147 1195 151
rect 1176 139 1180 143
rect 1288 102 1292 106
rect 1133 57 1137 61
rect 1149 59 1153 63
rect 1359 191 1363 195
rect 1494 195 1498 199
rect 1314 181 1318 185
rect 1344 183 1348 187
rect 1479 187 1483 191
rect 1541 193 1545 197
rect 1426 147 1430 151
rect 1411 139 1415 143
rect 1314 106 1318 110
rect 1302 65 1306 69
rect 1357 57 1361 61
rect 1385 57 1389 61
rect 1290 49 1294 53
rect 1342 49 1346 53
rect 1475 65 1479 69
rect 1459 49 1463 53
rect 1502 57 1506 61
rect 1578 377 1582 381
rect 1714 230 1718 234
rect 1699 222 1703 226
rect 1949 230 1953 234
rect 1934 222 1938 226
rect 1578 193 1582 197
rect 1570 185 1574 189
rect 1604 193 1608 197
rect 1647 191 1651 195
rect 1782 195 1786 199
rect 1604 181 1608 185
rect 1632 183 1636 187
rect 1767 187 1771 191
rect 1823 193 1827 197
rect 1714 147 1718 151
rect 1699 139 1703 143
rect 1811 102 1815 106
rect 1656 57 1660 61
rect 1672 59 1676 63
rect 1882 191 1886 195
rect 2017 195 2021 199
rect 1837 181 1841 185
rect 1867 183 1871 187
rect 2002 187 2006 191
rect 2064 193 2068 197
rect 1949 147 1953 151
rect 1934 139 1938 143
rect 1837 106 1841 110
rect 1825 65 1829 69
rect 1880 57 1884 61
rect 1908 57 1912 61
rect 1813 49 1817 53
rect 1865 49 1869 53
rect 1998 65 2002 69
rect 1982 49 1986 53
rect 2025 57 2029 61
<< ndcontact >>
rect -140 395 -136 399
rect -110 395 -106 399
rect -207 356 -203 360
rect -177 356 -173 360
rect -72 360 -68 364
rect -42 360 -38 364
rect -140 312 -136 316
rect -110 312 -106 316
rect 373 395 377 399
rect 403 395 407 399
rect 306 356 310 360
rect 336 356 340 360
rect 441 360 445 364
rect 471 360 475 364
rect 373 312 377 316
rect 403 312 407 316
rect 127 211 131 215
rect 157 211 161 215
rect 362 211 366 215
rect 60 172 64 176
rect 90 172 94 176
rect 195 176 199 180
rect 225 176 229 180
rect 127 128 131 132
rect 157 128 161 132
rect 41 38 45 42
rect 71 38 75 42
rect 83 38 87 42
rect 97 38 101 42
rect 392 211 396 215
rect 295 172 299 176
rect 325 172 329 176
rect 430 176 434 180
rect 460 176 464 180
rect 362 128 366 132
rect 392 128 396 132
rect 293 38 297 42
rect 323 38 327 42
rect 335 38 339 42
rect 349 38 353 42
rect 410 38 414 42
rect 424 38 428 42
rect 440 38 444 42
rect 452 38 456 42
rect 466 38 470 42
rect 879 395 883 399
rect 909 395 913 399
rect 812 356 816 360
rect 842 356 846 360
rect 947 360 951 364
rect 977 360 981 364
rect 879 312 883 316
rect 909 312 913 316
rect 650 211 654 215
rect 680 211 684 215
rect 885 211 889 215
rect 583 172 587 176
rect 613 172 617 176
rect 718 176 722 180
rect 748 176 752 180
rect 650 128 654 132
rect 680 128 684 132
rect 564 38 568 42
rect 594 38 598 42
rect 606 38 610 42
rect 620 38 624 42
rect 915 211 919 215
rect 818 172 822 176
rect 848 172 852 176
rect 953 176 957 180
rect 983 176 987 180
rect 885 128 889 132
rect 915 128 919 132
rect 816 38 820 42
rect 846 38 850 42
rect 858 38 862 42
rect 872 38 876 42
rect 933 38 937 42
rect 947 38 951 42
rect 963 38 967 42
rect 975 38 979 42
rect 989 38 993 42
rect 1403 395 1407 399
rect 1433 395 1437 399
rect 1336 356 1340 360
rect 1366 356 1370 360
rect 1471 360 1475 364
rect 1501 360 1505 364
rect 1403 312 1407 316
rect 1433 312 1437 316
rect 1173 211 1177 215
rect 1203 211 1207 215
rect 1408 211 1412 215
rect 1106 172 1110 176
rect 1136 172 1140 176
rect 1241 176 1245 180
rect 1271 176 1275 180
rect 1173 128 1177 132
rect 1203 128 1207 132
rect 1087 38 1091 42
rect 1117 38 1121 42
rect 1129 38 1133 42
rect 1143 38 1147 42
rect 1438 211 1442 215
rect 1341 172 1345 176
rect 1371 172 1375 176
rect 1476 176 1480 180
rect 1506 176 1510 180
rect 1408 128 1412 132
rect 1438 128 1442 132
rect 1339 38 1343 42
rect 1369 38 1373 42
rect 1381 38 1385 42
rect 1395 38 1399 42
rect 1456 38 1460 42
rect 1470 38 1474 42
rect 1486 38 1490 42
rect 1498 38 1502 42
rect 1512 38 1516 42
rect 1696 211 1700 215
rect 1726 211 1730 215
rect 1931 211 1935 215
rect 1629 172 1633 176
rect 1659 172 1663 176
rect 1764 176 1768 180
rect 1794 176 1798 180
rect 1696 128 1700 132
rect 1726 128 1730 132
rect 1610 38 1614 42
rect 1640 38 1644 42
rect 1652 38 1656 42
rect 1666 38 1670 42
rect 1961 211 1965 215
rect 1864 172 1868 176
rect 1894 172 1898 176
rect 1999 176 2003 180
rect 2029 176 2033 180
rect 1931 128 1935 132
rect 1961 128 1965 132
rect 1862 38 1866 42
rect 1892 38 1896 42
rect 1904 38 1908 42
rect 1918 38 1922 42
rect 1979 38 1983 42
rect 1993 38 1997 42
rect 2009 38 2013 42
rect 2021 38 2025 42
rect 2035 38 2039 42
<< pdcontact >>
rect -140 435 -136 439
rect -125 435 -121 439
rect -110 435 -106 439
rect -207 396 -203 400
rect -192 396 -188 400
rect -177 396 -173 400
rect -72 400 -68 404
rect -57 400 -53 404
rect -42 400 -38 404
rect -140 352 -136 356
rect -125 352 -121 356
rect -110 352 -106 356
rect 373 435 377 439
rect 388 435 392 439
rect 403 435 407 439
rect 306 396 310 400
rect 321 396 325 400
rect 336 396 340 400
rect 441 400 445 404
rect 456 400 460 404
rect 471 400 475 404
rect 373 352 377 356
rect 388 352 392 356
rect 403 352 407 356
rect 127 251 131 255
rect 142 251 146 255
rect 157 251 161 255
rect 362 251 366 255
rect 377 251 381 255
rect 392 251 396 255
rect 60 212 64 216
rect 75 212 79 216
rect 90 212 94 216
rect 195 216 199 220
rect 210 216 214 220
rect 225 216 229 220
rect 295 212 299 216
rect 310 212 314 216
rect 325 212 329 216
rect 127 168 131 172
rect 142 168 146 172
rect 157 168 161 172
rect 41 78 45 82
rect 56 78 60 82
rect 71 78 75 82
rect 83 78 87 82
rect 97 78 101 82
rect 430 216 434 220
rect 445 216 449 220
rect 460 216 464 220
rect 362 168 366 172
rect 377 168 381 172
rect 392 168 396 172
rect 293 78 297 82
rect 308 78 312 82
rect 323 78 327 82
rect 335 78 339 82
rect 349 78 353 82
rect 410 78 414 82
rect 440 78 444 82
rect 452 78 456 82
rect 466 78 470 82
rect 879 435 883 439
rect 894 435 898 439
rect 909 435 913 439
rect 812 396 816 400
rect 827 396 831 400
rect 842 396 846 400
rect 947 400 951 404
rect 962 400 966 404
rect 977 400 981 404
rect 879 352 883 356
rect 894 352 898 356
rect 909 352 913 356
rect 650 251 654 255
rect 665 251 669 255
rect 680 251 684 255
rect 885 251 889 255
rect 900 251 904 255
rect 915 251 919 255
rect 583 212 587 216
rect 598 212 602 216
rect 613 212 617 216
rect 718 216 722 220
rect 733 216 737 220
rect 748 216 752 220
rect 818 212 822 216
rect 833 212 837 216
rect 848 212 852 216
rect 650 168 654 172
rect 665 168 669 172
rect 680 168 684 172
rect 564 78 568 82
rect 579 78 583 82
rect 594 78 598 82
rect 606 78 610 82
rect 620 78 624 82
rect 953 216 957 220
rect 968 216 972 220
rect 983 216 987 220
rect 885 168 889 172
rect 900 168 904 172
rect 915 168 919 172
rect 816 78 820 82
rect 831 78 835 82
rect 846 78 850 82
rect 858 78 862 82
rect 872 78 876 82
rect 933 78 937 82
rect 963 78 967 82
rect 975 78 979 82
rect 989 78 993 82
rect 1403 435 1407 439
rect 1418 435 1422 439
rect 1433 435 1437 439
rect 1336 396 1340 400
rect 1351 396 1355 400
rect 1366 396 1370 400
rect 1471 400 1475 404
rect 1486 400 1490 404
rect 1501 400 1505 404
rect 1403 352 1407 356
rect 1418 352 1422 356
rect 1433 352 1437 356
rect 1173 251 1177 255
rect 1188 251 1192 255
rect 1203 251 1207 255
rect 1408 251 1412 255
rect 1423 251 1427 255
rect 1438 251 1442 255
rect 1106 212 1110 216
rect 1121 212 1125 216
rect 1136 212 1140 216
rect 1241 216 1245 220
rect 1256 216 1260 220
rect 1271 216 1275 220
rect 1341 212 1345 216
rect 1356 212 1360 216
rect 1371 212 1375 216
rect 1173 168 1177 172
rect 1188 168 1192 172
rect 1203 168 1207 172
rect 1087 78 1091 82
rect 1102 78 1106 82
rect 1117 78 1121 82
rect 1129 78 1133 82
rect 1143 78 1147 82
rect 1476 216 1480 220
rect 1491 216 1495 220
rect 1506 216 1510 220
rect 1408 168 1412 172
rect 1423 168 1427 172
rect 1438 168 1442 172
rect 1339 78 1343 82
rect 1354 78 1358 82
rect 1369 78 1373 82
rect 1381 78 1385 82
rect 1395 78 1399 82
rect 1456 78 1460 82
rect 1486 78 1490 82
rect 1498 78 1502 82
rect 1512 78 1516 82
rect 1696 251 1700 255
rect 1711 251 1715 255
rect 1726 251 1730 255
rect 1931 251 1935 255
rect 1946 251 1950 255
rect 1961 251 1965 255
rect 1629 212 1633 216
rect 1644 212 1648 216
rect 1659 212 1663 216
rect 1764 216 1768 220
rect 1779 216 1783 220
rect 1794 216 1798 220
rect 1864 212 1868 216
rect 1879 212 1883 216
rect 1894 212 1898 216
rect 1696 168 1700 172
rect 1711 168 1715 172
rect 1726 168 1730 172
rect 1610 78 1614 82
rect 1625 78 1629 82
rect 1640 78 1644 82
rect 1652 78 1656 82
rect 1666 78 1670 82
rect 1999 216 2003 220
rect 2014 216 2018 220
rect 2029 216 2033 220
rect 1931 168 1935 172
rect 1946 168 1950 172
rect 1961 168 1965 172
rect 1862 78 1866 82
rect 1877 78 1881 82
rect 1892 78 1896 82
rect 1904 78 1908 82
rect 1918 78 1922 82
rect 1979 78 1983 82
rect 2009 78 2013 82
rect 2021 78 2025 82
rect 2035 78 2039 82
<< nbccdiffcontact >>
rect 83 92 87 96
rect 335 92 339 96
rect 452 92 456 96
rect 606 92 610 96
rect 858 92 862 96
rect 975 92 979 96
rect 1129 92 1133 96
rect 1381 92 1385 96
rect 1498 92 1502 96
rect 1652 92 1656 96
rect 1904 92 1908 96
rect 2021 92 2025 96
<< m2contact >>
rect -172 447 -168 451
rect 341 447 345 451
rect 847 447 851 451
rect 1371 447 1375 451
rect -174 410 -170 414
rect -106 383 -102 387
rect -172 344 -168 348
rect -145 366 -141 370
rect 339 410 343 414
rect 407 383 411 387
rect -76 348 -72 352
rect 341 344 345 348
rect 368 366 372 370
rect 845 410 849 414
rect 913 383 917 387
rect 437 348 441 352
rect 847 344 851 348
rect 874 366 878 370
rect 1369 410 1373 414
rect 1437 383 1441 387
rect 943 348 947 352
rect 1371 344 1375 348
rect 1398 366 1402 370
rect 1467 348 1471 352
rect -162 302 -158 306
rect -102 302 -98 306
rect -78 302 -74 306
rect 351 302 355 306
rect -37 298 -33 302
rect 411 302 415 306
rect 435 302 439 306
rect 857 302 861 306
rect 917 302 921 306
rect 941 302 945 306
rect 1381 302 1385 306
rect 1441 302 1445 306
rect 1465 302 1469 306
rect 95 263 99 267
rect 330 263 334 267
rect 486 263 490 267
rect 618 263 622 267
rect 853 263 857 267
rect 1009 263 1013 267
rect 1141 263 1145 267
rect 1376 263 1380 267
rect 1532 263 1536 267
rect 1664 263 1668 267
rect 1899 263 1903 267
rect 2055 263 2059 267
rect 93 226 97 230
rect 161 199 165 203
rect 328 226 332 230
rect 95 160 99 164
rect 122 182 126 186
rect 396 199 400 203
rect 191 164 195 168
rect 330 160 334 164
rect 357 182 361 186
rect 616 226 620 230
rect 684 199 688 203
rect 851 226 855 230
rect 426 164 430 168
rect 618 160 622 164
rect 645 182 649 186
rect 919 199 923 203
rect 714 164 718 168
rect 853 160 857 164
rect 880 182 884 186
rect 1139 226 1143 230
rect 1207 199 1211 203
rect 1374 226 1378 230
rect 949 164 953 168
rect 1141 160 1145 164
rect 1168 182 1172 186
rect 1442 199 1446 203
rect 1237 164 1241 168
rect 1376 160 1380 164
rect 1403 182 1407 186
rect 1662 226 1666 230
rect 1730 199 1734 203
rect 1897 226 1901 230
rect 1472 164 1476 168
rect 1664 160 1668 164
rect 1691 182 1695 186
rect 1965 199 1969 203
rect 1760 164 1764 168
rect 1899 160 1903 164
rect 1926 182 1930 186
rect 1995 164 1999 168
rect 105 118 109 122
rect 165 118 169 122
rect 189 118 193 122
rect 340 118 344 122
rect 400 118 404 122
rect 424 118 428 122
rect 478 114 482 118
rect 628 118 632 122
rect 688 118 692 122
rect 712 118 716 122
rect 863 118 867 122
rect 923 118 927 122
rect 947 118 951 122
rect 1001 114 1005 118
rect 1151 118 1155 122
rect 1211 118 1215 122
rect 1235 118 1239 122
rect 1386 118 1390 122
rect 1446 118 1450 122
rect 1470 118 1474 122
rect 1524 114 1528 118
rect 1674 118 1678 122
rect 1734 118 1738 122
rect 1758 118 1762 122
rect 1909 118 1913 122
rect 1969 118 1973 122
rect 1993 118 1997 122
rect 2047 114 2051 118
rect 486 94 490 98
rect 1009 94 1013 98
rect 1532 94 1536 98
rect 2055 94 2059 98
rect -13 28 -9 32
rect 478 28 482 32
rect 1001 28 1005 32
rect 1524 28 1528 32
rect 2047 28 2051 32
<< psubstratepcontact >>
rect -135 383 -131 387
rect -114 383 -110 387
rect -202 344 -198 348
rect -181 344 -177 348
rect -67 348 -63 352
rect -46 348 -42 352
rect -135 300 -131 304
rect -114 300 -110 304
rect 378 383 382 387
rect 399 383 403 387
rect 311 344 315 348
rect 332 344 336 348
rect 446 348 450 352
rect 467 348 471 352
rect 378 300 382 304
rect 399 300 403 304
rect 132 199 136 203
rect 153 199 157 203
rect 65 160 69 164
rect 86 160 90 164
rect 200 164 204 168
rect 221 164 225 168
rect 132 116 136 120
rect 153 116 157 120
rect 46 26 50 30
rect 67 26 71 30
rect 83 26 87 30
rect 98 26 102 30
rect 367 199 371 203
rect 388 199 392 203
rect 300 160 304 164
rect 321 160 325 164
rect 435 164 439 168
rect 456 164 460 168
rect 367 116 371 120
rect 388 116 392 120
rect 298 26 302 30
rect 319 26 323 30
rect 335 26 339 30
rect 350 26 354 30
rect 415 26 419 30
rect 436 26 440 30
rect 452 26 456 30
rect 467 26 471 30
rect 884 383 888 387
rect 905 383 909 387
rect 817 344 821 348
rect 838 344 842 348
rect 952 348 956 352
rect 973 348 977 352
rect 884 300 888 304
rect 905 300 909 304
rect 655 199 659 203
rect 676 199 680 203
rect 588 160 592 164
rect 609 160 613 164
rect 723 164 727 168
rect 744 164 748 168
rect 655 116 659 120
rect 676 116 680 120
rect 569 26 573 30
rect 590 26 594 30
rect 606 26 610 30
rect 621 26 625 30
rect 890 199 894 203
rect 911 199 915 203
rect 823 160 827 164
rect 844 160 848 164
rect 958 164 962 168
rect 979 164 983 168
rect 890 116 894 120
rect 911 116 915 120
rect 821 26 825 30
rect 842 26 846 30
rect 858 26 862 30
rect 873 26 877 30
rect 938 26 942 30
rect 959 26 963 30
rect 975 26 979 30
rect 990 26 994 30
rect 1408 383 1412 387
rect 1429 383 1433 387
rect 1341 344 1345 348
rect 1362 344 1366 348
rect 1476 348 1480 352
rect 1497 348 1501 352
rect 1408 300 1412 304
rect 1429 300 1433 304
rect 1178 199 1182 203
rect 1199 199 1203 203
rect 1111 160 1115 164
rect 1132 160 1136 164
rect 1246 164 1250 168
rect 1267 164 1271 168
rect 1178 116 1182 120
rect 1199 116 1203 120
rect 1092 26 1096 30
rect 1113 26 1117 30
rect 1129 26 1133 30
rect 1144 26 1148 30
rect 1413 199 1417 203
rect 1434 199 1438 203
rect 1346 160 1350 164
rect 1367 160 1371 164
rect 1481 164 1485 168
rect 1502 164 1506 168
rect 1413 116 1417 120
rect 1434 116 1438 120
rect 1344 26 1348 30
rect 1365 26 1369 30
rect 1381 26 1385 30
rect 1396 26 1400 30
rect 1461 26 1465 30
rect 1482 26 1486 30
rect 1498 26 1502 30
rect 1513 26 1517 30
rect 1701 199 1705 203
rect 1722 199 1726 203
rect 1634 160 1638 164
rect 1655 160 1659 164
rect 1769 164 1773 168
rect 1790 164 1794 168
rect 1701 116 1705 120
rect 1722 116 1726 120
rect 1615 26 1619 30
rect 1636 26 1640 30
rect 1652 26 1656 30
rect 1667 26 1671 30
rect 1936 199 1940 203
rect 1957 199 1961 203
rect 1869 160 1873 164
rect 1890 160 1894 164
rect 2004 164 2008 168
rect 2025 164 2029 168
rect 1936 116 1940 120
rect 1957 116 1961 120
rect 1867 26 1871 30
rect 1888 26 1892 30
rect 1904 26 1908 30
rect 1919 26 1923 30
rect 1984 26 1988 30
rect 2005 26 2009 30
rect 2021 26 2025 30
rect 2036 26 2040 30
<< nsubstratencontact >>
rect -135 449 -131 453
rect -116 449 -112 453
rect -202 410 -198 414
rect -183 410 -179 414
rect -67 414 -63 418
rect -48 414 -44 418
rect -135 366 -131 370
rect -116 366 -112 370
rect 378 449 382 453
rect 397 449 401 453
rect 311 410 315 414
rect 330 410 334 414
rect 446 414 450 418
rect 465 414 469 418
rect 378 366 382 370
rect 397 366 401 370
rect 132 265 136 269
rect 151 265 155 269
rect 367 265 371 269
rect 386 265 390 269
rect 65 226 69 230
rect 84 226 88 230
rect 200 230 204 234
rect 219 230 223 234
rect 300 226 304 230
rect 319 226 323 230
rect 435 230 439 234
rect 454 230 458 234
rect 132 182 136 186
rect 151 182 155 186
rect 46 92 50 96
rect 65 92 69 96
rect 97 92 101 96
rect 367 182 371 186
rect 386 182 390 186
rect 298 92 302 96
rect 317 92 321 96
rect 349 92 353 96
rect 415 92 419 96
rect 434 92 438 96
rect 466 92 470 96
rect 884 449 888 453
rect 903 449 907 453
rect 817 410 821 414
rect 836 410 840 414
rect 952 414 956 418
rect 971 414 975 418
rect 884 366 888 370
rect 903 366 907 370
rect 655 265 659 269
rect 674 265 678 269
rect 890 265 894 269
rect 909 265 913 269
rect 588 226 592 230
rect 607 226 611 230
rect 723 230 727 234
rect 742 230 746 234
rect 823 226 827 230
rect 842 226 846 230
rect 958 230 962 234
rect 977 230 981 234
rect 655 182 659 186
rect 674 182 678 186
rect 569 92 573 96
rect 588 92 592 96
rect 620 92 624 96
rect 890 182 894 186
rect 909 182 913 186
rect 821 92 825 96
rect 840 92 844 96
rect 872 92 876 96
rect 938 92 942 96
rect 957 92 961 96
rect 989 92 993 96
rect 1408 449 1412 453
rect 1427 449 1431 453
rect 1341 410 1345 414
rect 1360 410 1364 414
rect 1476 414 1480 418
rect 1495 414 1499 418
rect 1408 366 1412 370
rect 1427 366 1431 370
rect 1178 265 1182 269
rect 1197 265 1201 269
rect 1413 265 1417 269
rect 1432 265 1436 269
rect 1111 226 1115 230
rect 1130 226 1134 230
rect 1246 230 1250 234
rect 1265 230 1269 234
rect 1346 226 1350 230
rect 1365 226 1369 230
rect 1481 230 1485 234
rect 1500 230 1504 234
rect 1178 182 1182 186
rect 1197 182 1201 186
rect 1092 92 1096 96
rect 1111 92 1115 96
rect 1143 92 1147 96
rect 1413 182 1417 186
rect 1432 182 1436 186
rect 1344 92 1348 96
rect 1363 92 1367 96
rect 1395 92 1399 96
rect 1461 92 1465 96
rect 1480 92 1484 96
rect 1512 92 1516 96
rect 1701 265 1705 269
rect 1720 265 1724 269
rect 1936 265 1940 269
rect 1955 265 1959 269
rect 1634 226 1638 230
rect 1653 226 1657 230
rect 1769 230 1773 234
rect 1788 230 1792 234
rect 1869 226 1873 230
rect 1888 226 1892 230
rect 2004 230 2008 234
rect 2023 230 2027 234
rect 1701 182 1705 186
rect 1720 182 1724 186
rect 1615 92 1619 96
rect 1634 92 1638 96
rect 1666 92 1670 96
rect 1936 182 1940 186
rect 1955 182 1959 186
rect 1867 92 1871 96
rect 1886 92 1890 96
rect 1918 92 1922 96
rect 1984 92 1988 96
rect 2003 92 2007 96
rect 2035 92 2039 96
<< labels >>
rlabel metal1 560 266 560 266 1 Vdd
rlabel metal1 552 28 552 28 1 gnd
rlabel polysilicon 3 278 3 278 5 a0
rlabel polysilicon 526 277 526 277 5 a1
rlabel polysilicon 1049 276 1049 276 5 a2
rlabel polysilicon 1572 276 1572 276 5 a3
rlabel metal1 2077 61 2077 61 7 Carry
rlabel polysilicon 2066 13 2066 13 1 s3
rlabel polysilicon 1543 14 1543 14 1 s2
rlabel polysilicon 1020 14 1020 14 1 s1
rlabel polysilicon 497 14 497 14 1 s0
rlabel polysilicon -276 467 -276 467 4 b0
rlabel polysilicon 282 467 282 467 5 b1
rlabel polysilicon 787 466 787 466 5 b2
rlabel polysilicon 1311 465 1311 465 5 b3
rlabel metal1 -242 285 -242 285 1 ctrl
<< end >>
