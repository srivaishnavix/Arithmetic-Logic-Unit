* SPICE3 file created from ANDGATE.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'


.option scale=1u

M1000 Vout a_15_50# Vdd w_0_48# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1001 Vout a_15_50# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1002 a_15_50# Va Vdd w_0_48# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1003 Vdd Vb a_15_50# w_0_48# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1004 a_15_10# Va gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1005 a_15_50# Vb a_15_10# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
C0 gnd 0 11.656f 
C1 Vout 0 6.392f 
C2 a_15_50# 0 21.108f 
C3 Vb 0 18.154f 
C4 Va 0 14.394f 
C5 Vdd 0 13.16f 



Va Va gnd 0
Vb Vb gnd 1


.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(Va) v(Vb)+2 v(Vout)+4 
.end
.endc