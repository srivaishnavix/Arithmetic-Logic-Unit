magic
tech scmos
timestamp 1700600272
<< nwell >>
rect 91 234 133 246
rect 305 238 347 250
rect 598 233 640 245
rect 812 237 854 249
rect 1108 233 1150 245
rect 1322 237 1364 249
rect 1647 233 1689 245
rect 1861 237 1903 249
rect 24 195 66 207
rect 159 199 201 211
rect 238 199 280 211
rect 373 203 415 215
rect 531 194 573 206
rect 666 198 708 210
rect 745 198 787 210
rect 880 202 922 214
rect 1041 194 1083 206
rect 1176 198 1218 210
rect 1255 198 1297 210
rect 1390 202 1432 214
rect 1580 194 1622 206
rect 1715 198 1757 210
rect 1794 198 1836 210
rect 1929 202 1971 214
rect 91 151 133 163
rect 305 155 347 167
rect 598 150 640 162
rect 812 154 854 166
rect 1108 150 1150 162
rect 1322 154 1364 166
rect 1647 150 1689 162
rect 1861 154 1903 166
rect 18 51 86 63
rect 240 51 308 63
rect 352 51 420 63
rect 525 50 593 62
rect 747 50 815 62
rect 859 50 927 62
rect 1035 50 1103 62
rect 1257 50 1325 62
rect 1369 50 1437 62
rect 1574 50 1642 62
rect 1796 50 1864 62
rect 1908 50 1976 62
<< polysilicon >>
rect 317 248 320 252
rect 332 248 335 252
rect 103 244 106 248
rect 118 244 121 248
rect 824 247 827 251
rect 839 247 842 251
rect 1334 247 1337 251
rect 1349 247 1352 251
rect 1873 247 1876 251
rect 1888 247 1891 251
rect 610 243 613 247
rect 625 243 628 247
rect 103 213 106 236
rect 118 221 121 236
rect 117 217 121 221
rect 317 217 320 240
rect 332 225 335 240
rect 1120 243 1123 247
rect 1135 243 1138 247
rect 331 221 335 225
rect 102 209 106 213
rect 36 205 39 209
rect 51 205 54 209
rect 103 204 106 209
rect 118 204 121 217
rect 316 213 320 217
rect 171 209 174 213
rect 186 209 189 213
rect 250 209 253 213
rect 265 209 268 213
rect -5 30 -1 168
rect 8 46 12 177
rect 36 174 39 197
rect 51 182 54 197
rect 317 208 320 213
rect 332 208 335 221
rect 385 213 388 217
rect 400 213 403 217
rect 103 194 106 196
rect 118 194 121 196
rect 50 178 54 182
rect 171 178 174 201
rect 186 186 189 201
rect 185 182 189 186
rect 35 170 39 174
rect 36 165 39 170
rect 51 165 54 178
rect 170 174 174 178
rect 171 169 174 174
rect 186 169 189 182
rect 103 161 106 165
rect 118 161 121 165
rect 36 155 39 157
rect 51 155 54 157
rect 171 159 174 161
rect 186 159 189 161
rect 103 130 106 153
rect 118 138 121 153
rect 117 134 121 138
rect 102 126 106 130
rect 103 121 106 126
rect 118 121 121 134
rect 103 111 106 113
rect 118 111 121 113
rect 30 61 33 65
rect 45 61 48 65
rect 72 61 74 65
rect 8 42 16 46
rect 30 30 33 53
rect 45 38 48 53
rect 44 34 48 38
rect -5 26 16 30
rect 29 26 33 30
rect 30 21 33 26
rect 45 21 48 34
rect 72 21 74 53
rect 88 36 121 40
rect 30 11 33 13
rect 45 11 48 13
rect 72 11 74 13
rect 117 1 121 36
rect 205 30 209 180
rect 250 178 253 201
rect 265 186 268 201
rect 610 212 613 235
rect 625 220 628 235
rect 624 216 628 220
rect 824 216 827 239
rect 839 224 842 239
rect 1659 243 1662 247
rect 1674 243 1677 247
rect 838 220 842 224
rect 609 208 613 212
rect 317 198 320 200
rect 332 198 335 200
rect 264 182 268 186
rect 385 182 388 205
rect 400 190 403 205
rect 543 204 546 208
rect 558 204 561 208
rect 610 203 613 208
rect 625 203 628 216
rect 823 212 827 216
rect 678 208 681 212
rect 693 208 696 212
rect 757 208 760 212
rect 772 208 775 212
rect 399 186 403 190
rect 444 186 461 190
rect 249 174 253 178
rect 250 169 253 174
rect 265 169 268 182
rect 384 178 388 182
rect 385 173 388 178
rect 400 173 403 186
rect 317 165 320 169
rect 332 165 335 169
rect 250 159 253 161
rect 265 159 268 161
rect 385 163 388 165
rect 400 163 403 165
rect 317 134 320 157
rect 332 142 335 157
rect 331 138 335 142
rect 316 130 320 134
rect 317 125 320 130
rect 332 125 335 138
rect 317 115 320 117
rect 332 115 335 117
rect 217 46 221 93
rect 252 61 255 65
rect 267 61 270 65
rect 294 61 296 65
rect 364 61 367 65
rect 379 61 382 65
rect 406 61 408 65
rect 217 42 238 46
rect 252 30 255 53
rect 267 38 270 53
rect 266 34 270 38
rect 205 26 237 30
rect 251 26 255 30
rect 252 21 255 26
rect 267 21 270 34
rect 294 21 296 53
rect 345 42 350 46
rect 345 40 349 42
rect 311 36 349 40
rect 364 30 367 53
rect 348 29 350 30
rect 323 26 350 29
rect 363 26 367 30
rect 323 25 354 26
rect 252 11 255 13
rect 267 11 270 13
rect 294 11 296 13
rect 323 1 327 25
rect 364 21 367 26
rect 379 21 382 53
rect 406 21 408 53
rect 364 11 367 13
rect 379 11 382 13
rect 406 11 408 13
rect 117 -3 327 1
rect 457 -77 461 186
rect 502 29 506 167
rect 515 45 519 176
rect 543 173 546 196
rect 558 181 561 196
rect 824 207 827 212
rect 839 207 842 220
rect 892 212 895 216
rect 907 212 910 216
rect 1120 212 1123 235
rect 1135 220 1138 235
rect 1134 216 1138 220
rect 1334 216 1337 239
rect 1349 224 1352 239
rect 1348 220 1352 224
rect 610 193 613 195
rect 625 193 628 195
rect 557 177 561 181
rect 678 177 681 200
rect 693 185 696 200
rect 692 181 696 185
rect 542 169 546 173
rect 543 164 546 169
rect 558 164 561 177
rect 677 173 681 177
rect 678 168 681 173
rect 693 168 696 181
rect 610 160 613 164
rect 625 160 628 164
rect 543 154 546 156
rect 558 154 561 156
rect 678 158 681 160
rect 693 158 696 160
rect 610 129 613 152
rect 625 137 628 152
rect 624 133 628 137
rect 609 125 613 129
rect 610 120 613 125
rect 625 120 628 133
rect 610 110 613 112
rect 625 110 628 112
rect 537 60 540 64
rect 552 60 555 64
rect 579 60 581 64
rect 515 41 523 45
rect 537 29 540 52
rect 552 37 555 52
rect 551 33 555 37
rect 502 25 523 29
rect 536 25 540 29
rect 537 20 540 25
rect 552 20 555 33
rect 579 20 581 52
rect 595 35 628 39
rect 537 10 540 12
rect 552 10 555 12
rect 579 10 581 12
rect 624 0 628 35
rect 712 29 716 179
rect 757 177 760 200
rect 772 185 775 200
rect 1119 208 1123 212
rect 1053 204 1056 208
rect 1068 204 1071 208
rect 824 197 827 199
rect 839 197 842 199
rect 771 181 775 185
rect 892 181 895 204
rect 907 189 910 204
rect 1120 203 1123 208
rect 1135 203 1138 216
rect 1333 212 1337 216
rect 1188 208 1191 212
rect 1203 208 1206 212
rect 1267 208 1270 212
rect 1282 208 1285 212
rect 906 185 910 189
rect 951 185 972 189
rect 756 173 760 177
rect 757 168 760 173
rect 772 168 775 181
rect 891 177 895 181
rect 892 172 895 177
rect 907 172 910 185
rect 824 164 827 168
rect 839 164 842 168
rect 757 158 760 160
rect 772 158 775 160
rect 892 162 895 164
rect 907 162 910 164
rect 824 133 827 156
rect 839 141 842 156
rect 838 137 842 141
rect 823 129 827 133
rect 824 124 827 129
rect 839 124 842 137
rect 824 114 827 116
rect 839 114 842 116
rect 724 45 728 92
rect 759 60 762 64
rect 774 60 777 64
rect 801 60 803 64
rect 871 60 874 64
rect 886 60 889 64
rect 913 60 915 64
rect 724 41 745 45
rect 759 29 762 52
rect 774 37 777 52
rect 773 33 777 37
rect 712 25 744 29
rect 758 25 762 29
rect 759 20 762 25
rect 774 20 777 33
rect 801 20 803 52
rect 852 41 857 45
rect 852 39 856 41
rect 818 35 856 39
rect 871 29 874 52
rect 855 28 857 29
rect 830 25 857 28
rect 870 25 874 29
rect 830 24 861 25
rect 759 10 762 12
rect 774 10 777 12
rect 801 10 803 12
rect 830 0 834 24
rect 871 20 874 25
rect 886 20 889 52
rect 913 20 915 52
rect 871 10 874 12
rect 886 10 889 12
rect 913 10 915 12
rect 624 -4 834 0
rect 968 -78 972 185
rect 1012 29 1016 167
rect 1025 45 1029 176
rect 1053 173 1056 196
rect 1068 181 1071 196
rect 1334 207 1337 212
rect 1349 207 1352 220
rect 1402 212 1405 216
rect 1417 212 1420 216
rect 1659 212 1662 235
rect 1674 220 1677 235
rect 1673 216 1677 220
rect 1873 216 1876 239
rect 1888 224 1891 239
rect 1887 220 1891 224
rect 1120 193 1123 195
rect 1135 193 1138 195
rect 1067 177 1071 181
rect 1188 177 1191 200
rect 1203 185 1206 200
rect 1202 181 1206 185
rect 1052 169 1056 173
rect 1053 164 1056 169
rect 1068 164 1071 177
rect 1187 173 1191 177
rect 1188 168 1191 173
rect 1203 168 1206 181
rect 1120 160 1123 164
rect 1135 160 1138 164
rect 1053 154 1056 156
rect 1068 154 1071 156
rect 1188 158 1191 160
rect 1203 158 1206 160
rect 1120 129 1123 152
rect 1135 137 1138 152
rect 1134 133 1138 137
rect 1119 125 1123 129
rect 1120 120 1123 125
rect 1135 120 1138 133
rect 1120 110 1123 112
rect 1135 110 1138 112
rect 1047 60 1050 64
rect 1062 60 1065 64
rect 1089 60 1091 64
rect 1025 41 1033 45
rect 1047 29 1050 52
rect 1062 37 1065 52
rect 1061 33 1065 37
rect 1012 25 1033 29
rect 1046 25 1050 29
rect 1047 20 1050 25
rect 1062 20 1065 33
rect 1089 20 1091 52
rect 1105 35 1138 39
rect 1047 10 1050 12
rect 1062 10 1065 12
rect 1089 10 1091 12
rect 1134 0 1138 35
rect 1222 29 1226 179
rect 1267 177 1270 200
rect 1282 185 1285 200
rect 1658 208 1662 212
rect 1592 204 1595 208
rect 1607 204 1610 208
rect 1334 197 1337 199
rect 1349 197 1352 199
rect 1281 181 1285 185
rect 1402 181 1405 204
rect 1417 189 1420 204
rect 1659 203 1662 208
rect 1674 203 1677 216
rect 1872 212 1876 216
rect 1727 208 1730 212
rect 1742 208 1745 212
rect 1806 208 1809 212
rect 1821 208 1824 212
rect 1416 185 1420 189
rect 1461 185 1493 189
rect 1266 173 1270 177
rect 1267 168 1270 173
rect 1282 168 1285 181
rect 1401 177 1405 181
rect 1402 172 1405 177
rect 1417 172 1420 185
rect 1334 164 1337 168
rect 1349 164 1352 168
rect 1267 158 1270 160
rect 1282 158 1285 160
rect 1402 162 1405 164
rect 1417 162 1420 164
rect 1334 133 1337 156
rect 1349 141 1352 156
rect 1348 137 1352 141
rect 1333 129 1337 133
rect 1334 124 1337 129
rect 1349 124 1352 137
rect 1334 114 1337 116
rect 1349 114 1352 116
rect 1234 45 1238 92
rect 1269 60 1272 64
rect 1284 60 1287 64
rect 1311 60 1313 64
rect 1381 60 1384 64
rect 1396 60 1399 64
rect 1423 60 1425 64
rect 1234 41 1255 45
rect 1269 29 1272 52
rect 1284 37 1287 52
rect 1283 33 1287 37
rect 1222 25 1254 29
rect 1268 25 1272 29
rect 1269 20 1272 25
rect 1284 20 1287 33
rect 1311 20 1313 52
rect 1362 41 1367 45
rect 1362 39 1366 41
rect 1328 35 1366 39
rect 1381 29 1384 52
rect 1365 28 1367 29
rect 1340 25 1367 28
rect 1380 25 1384 29
rect 1340 24 1371 25
rect 1269 10 1272 12
rect 1284 10 1287 12
rect 1311 10 1313 12
rect 1340 0 1344 24
rect 1381 20 1384 25
rect 1396 20 1399 52
rect 1423 20 1425 52
rect 1381 10 1384 12
rect 1396 10 1399 12
rect 1423 10 1425 12
rect 1134 -4 1344 0
rect 1489 -78 1493 185
rect 1551 29 1555 167
rect 1564 45 1568 176
rect 1592 173 1595 196
rect 1607 181 1610 196
rect 1873 207 1876 212
rect 1888 207 1891 220
rect 1941 212 1944 216
rect 1956 212 1959 216
rect 1659 193 1662 195
rect 1674 193 1677 195
rect 1606 177 1610 181
rect 1727 177 1730 200
rect 1742 185 1745 200
rect 1741 181 1745 185
rect 1591 169 1595 173
rect 1592 164 1595 169
rect 1607 164 1610 177
rect 1726 173 1730 177
rect 1727 168 1730 173
rect 1742 168 1745 181
rect 1659 160 1662 164
rect 1674 160 1677 164
rect 1592 154 1595 156
rect 1607 154 1610 156
rect 1727 158 1730 160
rect 1742 158 1745 160
rect 1659 129 1662 152
rect 1674 137 1677 152
rect 1673 133 1677 137
rect 1658 125 1662 129
rect 1659 120 1662 125
rect 1674 120 1677 133
rect 1659 110 1662 112
rect 1674 110 1677 112
rect 1586 60 1589 64
rect 1601 60 1604 64
rect 1628 60 1630 64
rect 1564 41 1572 45
rect 1586 29 1589 52
rect 1601 37 1604 52
rect 1600 33 1604 37
rect 1551 25 1572 29
rect 1585 25 1589 29
rect 1586 20 1589 25
rect 1601 20 1604 33
rect 1628 20 1630 52
rect 1644 35 1677 39
rect 1586 10 1589 12
rect 1601 10 1604 12
rect 1628 10 1630 12
rect 1673 0 1677 35
rect 1761 29 1765 179
rect 1806 177 1809 200
rect 1821 185 1824 200
rect 1873 197 1876 199
rect 1888 197 1891 199
rect 1820 181 1824 185
rect 1941 181 1944 204
rect 1956 189 1959 204
rect 1955 185 1959 189
rect 2000 185 2070 189
rect 1805 173 1809 177
rect 1806 168 1809 173
rect 1821 168 1824 181
rect 1940 177 1944 181
rect 1941 172 1944 177
rect 1956 172 1959 185
rect 1873 164 1876 168
rect 1888 164 1891 168
rect 2002 171 2037 175
rect 1806 158 1809 160
rect 1821 158 1824 160
rect 1941 162 1944 164
rect 1956 162 1959 164
rect 1873 133 1876 156
rect 1888 141 1891 156
rect 1887 137 1891 141
rect 1872 129 1876 133
rect 1873 124 1876 129
rect 1888 124 1891 137
rect 1873 114 1876 116
rect 1888 114 1891 116
rect 1773 45 1777 92
rect 1808 60 1811 64
rect 1823 60 1826 64
rect 1850 60 1852 64
rect 1920 60 1923 64
rect 1935 60 1938 64
rect 1962 60 1964 64
rect 1773 41 1794 45
rect 1808 29 1811 52
rect 1823 37 1826 52
rect 1822 33 1826 37
rect 1761 25 1793 29
rect 1807 25 1811 29
rect 1808 20 1811 25
rect 1823 20 1826 33
rect 1850 20 1852 52
rect 1901 41 1906 45
rect 1901 39 1905 41
rect 1867 35 1905 39
rect 1920 29 1923 52
rect 1904 28 1908 29
rect 1879 25 1908 28
rect 1919 25 1923 29
rect 1879 24 1910 25
rect 1808 10 1811 12
rect 1823 10 1826 12
rect 1850 10 1852 12
rect 1879 0 1883 24
rect 1920 20 1923 25
rect 1935 20 1938 52
rect 1962 20 1964 52
rect 1920 10 1923 12
rect 1935 10 1938 12
rect 1962 10 1964 12
rect 1673 -4 1883 0
rect 2033 -80 2037 171
rect 2066 -79 2070 185
<< ndiffusion >>
rect 93 202 103 204
rect 93 198 95 202
rect 99 198 103 202
rect 93 196 103 198
rect 106 196 118 204
rect 121 202 131 204
rect 121 198 125 202
rect 129 198 131 202
rect 307 206 317 208
rect 307 202 309 206
rect 313 202 317 206
rect 121 196 131 198
rect 161 167 171 169
rect 26 163 36 165
rect 26 159 28 163
rect 32 159 36 163
rect 26 157 36 159
rect 39 157 51 165
rect 54 163 64 165
rect 54 159 58 163
rect 62 159 64 163
rect 161 163 163 167
rect 167 163 171 167
rect 161 161 171 163
rect 174 161 186 169
rect 189 167 199 169
rect 189 163 193 167
rect 197 163 199 167
rect 189 161 199 163
rect 54 157 64 159
rect 93 119 103 121
rect 93 115 95 119
rect 99 115 103 119
rect 93 113 103 115
rect 106 113 118 121
rect 121 119 131 121
rect 121 115 125 119
rect 129 115 131 119
rect 121 113 131 115
rect 20 19 30 21
rect 20 15 22 19
rect 26 15 30 19
rect 20 13 30 15
rect 33 13 45 21
rect 48 19 58 21
rect 48 15 52 19
rect 56 15 58 19
rect 48 13 58 15
rect 62 19 72 21
rect 62 15 64 19
rect 68 15 72 19
rect 62 13 72 15
rect 74 19 84 21
rect 74 15 78 19
rect 82 15 84 19
rect 74 13 84 15
rect 307 200 317 202
rect 320 200 332 208
rect 335 206 345 208
rect 335 202 339 206
rect 343 202 345 206
rect 335 200 345 202
rect 600 201 610 203
rect 600 197 602 201
rect 606 197 610 201
rect 375 171 385 173
rect 240 167 250 169
rect 240 163 242 167
rect 246 163 250 167
rect 240 161 250 163
rect 253 161 265 169
rect 268 167 278 169
rect 268 163 272 167
rect 276 163 278 167
rect 375 167 377 171
rect 381 167 385 171
rect 375 165 385 167
rect 388 165 400 173
rect 403 171 413 173
rect 403 167 407 171
rect 411 167 413 171
rect 403 165 413 167
rect 268 161 278 163
rect 307 123 317 125
rect 307 119 309 123
rect 313 119 317 123
rect 307 117 317 119
rect 320 117 332 125
rect 335 123 345 125
rect 335 119 339 123
rect 343 119 345 123
rect 335 117 345 119
rect 242 19 252 21
rect 242 15 244 19
rect 248 15 252 19
rect 242 13 252 15
rect 255 13 267 21
rect 270 19 280 21
rect 270 15 274 19
rect 278 15 280 19
rect 270 13 280 15
rect 284 19 294 21
rect 284 15 286 19
rect 290 15 294 19
rect 284 13 294 15
rect 296 19 306 21
rect 296 15 300 19
rect 304 15 306 19
rect 296 13 306 15
rect 354 19 364 21
rect 354 15 356 19
rect 360 15 364 19
rect 354 13 364 15
rect 367 19 379 21
rect 367 15 370 19
rect 374 15 379 19
rect 367 13 379 15
rect 382 19 392 21
rect 382 15 386 19
rect 390 15 392 19
rect 382 13 392 15
rect 396 19 406 21
rect 396 15 398 19
rect 402 15 406 19
rect 396 13 406 15
rect 408 19 418 21
rect 408 15 412 19
rect 416 15 418 19
rect 408 13 418 15
rect 600 195 610 197
rect 613 195 625 203
rect 628 201 638 203
rect 628 197 632 201
rect 636 197 638 201
rect 814 205 824 207
rect 814 201 816 205
rect 820 201 824 205
rect 628 195 638 197
rect 668 166 678 168
rect 533 162 543 164
rect 533 158 535 162
rect 539 158 543 162
rect 533 156 543 158
rect 546 156 558 164
rect 561 162 571 164
rect 561 158 565 162
rect 569 158 571 162
rect 668 162 670 166
rect 674 162 678 166
rect 668 160 678 162
rect 681 160 693 168
rect 696 166 706 168
rect 696 162 700 166
rect 704 162 706 166
rect 696 160 706 162
rect 561 156 571 158
rect 600 118 610 120
rect 600 114 602 118
rect 606 114 610 118
rect 600 112 610 114
rect 613 112 625 120
rect 628 118 638 120
rect 628 114 632 118
rect 636 114 638 118
rect 628 112 638 114
rect 527 18 537 20
rect 527 14 529 18
rect 533 14 537 18
rect 527 12 537 14
rect 540 12 552 20
rect 555 18 565 20
rect 555 14 559 18
rect 563 14 565 18
rect 555 12 565 14
rect 569 18 579 20
rect 569 14 571 18
rect 575 14 579 18
rect 569 12 579 14
rect 581 18 591 20
rect 581 14 585 18
rect 589 14 591 18
rect 581 12 591 14
rect 814 199 824 201
rect 827 199 839 207
rect 842 205 852 207
rect 842 201 846 205
rect 850 201 852 205
rect 842 199 852 201
rect 1110 201 1120 203
rect 1110 197 1112 201
rect 1116 197 1120 201
rect 882 170 892 172
rect 747 166 757 168
rect 747 162 749 166
rect 753 162 757 166
rect 747 160 757 162
rect 760 160 772 168
rect 775 166 785 168
rect 775 162 779 166
rect 783 162 785 166
rect 882 166 884 170
rect 888 166 892 170
rect 882 164 892 166
rect 895 164 907 172
rect 910 170 920 172
rect 910 166 914 170
rect 918 166 920 170
rect 910 164 920 166
rect 775 160 785 162
rect 814 122 824 124
rect 814 118 816 122
rect 820 118 824 122
rect 814 116 824 118
rect 827 116 839 124
rect 842 122 852 124
rect 842 118 846 122
rect 850 118 852 122
rect 842 116 852 118
rect 749 18 759 20
rect 749 14 751 18
rect 755 14 759 18
rect 749 12 759 14
rect 762 12 774 20
rect 777 18 787 20
rect 777 14 781 18
rect 785 14 787 18
rect 777 12 787 14
rect 791 18 801 20
rect 791 14 793 18
rect 797 14 801 18
rect 791 12 801 14
rect 803 18 813 20
rect 803 14 807 18
rect 811 14 813 18
rect 803 12 813 14
rect 861 18 871 20
rect 861 14 863 18
rect 867 14 871 18
rect 861 12 871 14
rect 874 18 886 20
rect 874 14 877 18
rect 881 14 886 18
rect 874 12 886 14
rect 889 18 899 20
rect 889 14 893 18
rect 897 14 899 18
rect 889 12 899 14
rect 903 18 913 20
rect 903 14 905 18
rect 909 14 913 18
rect 903 12 913 14
rect 915 18 925 20
rect 915 14 919 18
rect 923 14 925 18
rect 915 12 925 14
rect 1110 195 1120 197
rect 1123 195 1135 203
rect 1138 201 1148 203
rect 1138 197 1142 201
rect 1146 197 1148 201
rect 1324 205 1334 207
rect 1324 201 1326 205
rect 1330 201 1334 205
rect 1138 195 1148 197
rect 1178 166 1188 168
rect 1043 162 1053 164
rect 1043 158 1045 162
rect 1049 158 1053 162
rect 1043 156 1053 158
rect 1056 156 1068 164
rect 1071 162 1081 164
rect 1071 158 1075 162
rect 1079 158 1081 162
rect 1178 162 1180 166
rect 1184 162 1188 166
rect 1178 160 1188 162
rect 1191 160 1203 168
rect 1206 166 1216 168
rect 1206 162 1210 166
rect 1214 162 1216 166
rect 1206 160 1216 162
rect 1071 156 1081 158
rect 1110 118 1120 120
rect 1110 114 1112 118
rect 1116 114 1120 118
rect 1110 112 1120 114
rect 1123 112 1135 120
rect 1138 118 1148 120
rect 1138 114 1142 118
rect 1146 114 1148 118
rect 1138 112 1148 114
rect 1037 18 1047 20
rect 1037 14 1039 18
rect 1043 14 1047 18
rect 1037 12 1047 14
rect 1050 12 1062 20
rect 1065 18 1075 20
rect 1065 14 1069 18
rect 1073 14 1075 18
rect 1065 12 1075 14
rect 1079 18 1089 20
rect 1079 14 1081 18
rect 1085 14 1089 18
rect 1079 12 1089 14
rect 1091 18 1101 20
rect 1091 14 1095 18
rect 1099 14 1101 18
rect 1091 12 1101 14
rect 1324 199 1334 201
rect 1337 199 1349 207
rect 1352 205 1362 207
rect 1352 201 1356 205
rect 1360 201 1362 205
rect 1352 199 1362 201
rect 1649 201 1659 203
rect 1649 197 1651 201
rect 1655 197 1659 201
rect 1392 170 1402 172
rect 1257 166 1267 168
rect 1257 162 1259 166
rect 1263 162 1267 166
rect 1257 160 1267 162
rect 1270 160 1282 168
rect 1285 166 1295 168
rect 1285 162 1289 166
rect 1293 162 1295 166
rect 1392 166 1394 170
rect 1398 166 1402 170
rect 1392 164 1402 166
rect 1405 164 1417 172
rect 1420 170 1430 172
rect 1420 166 1424 170
rect 1428 166 1430 170
rect 1420 164 1430 166
rect 1285 160 1295 162
rect 1324 122 1334 124
rect 1324 118 1326 122
rect 1330 118 1334 122
rect 1324 116 1334 118
rect 1337 116 1349 124
rect 1352 122 1362 124
rect 1352 118 1356 122
rect 1360 118 1362 122
rect 1352 116 1362 118
rect 1259 18 1269 20
rect 1259 14 1261 18
rect 1265 14 1269 18
rect 1259 12 1269 14
rect 1272 12 1284 20
rect 1287 18 1297 20
rect 1287 14 1291 18
rect 1295 14 1297 18
rect 1287 12 1297 14
rect 1301 18 1311 20
rect 1301 14 1303 18
rect 1307 14 1311 18
rect 1301 12 1311 14
rect 1313 18 1323 20
rect 1313 14 1317 18
rect 1321 14 1323 18
rect 1313 12 1323 14
rect 1371 18 1381 20
rect 1371 14 1373 18
rect 1377 14 1381 18
rect 1371 12 1381 14
rect 1384 18 1396 20
rect 1384 14 1387 18
rect 1391 14 1396 18
rect 1384 12 1396 14
rect 1399 18 1409 20
rect 1399 14 1403 18
rect 1407 14 1409 18
rect 1399 12 1409 14
rect 1413 18 1423 20
rect 1413 14 1415 18
rect 1419 14 1423 18
rect 1413 12 1423 14
rect 1425 18 1435 20
rect 1425 14 1429 18
rect 1433 14 1435 18
rect 1425 12 1435 14
rect 1649 195 1659 197
rect 1662 195 1674 203
rect 1677 201 1687 203
rect 1677 197 1681 201
rect 1685 197 1687 201
rect 1863 205 1873 207
rect 1863 201 1865 205
rect 1869 201 1873 205
rect 1677 195 1687 197
rect 1717 166 1727 168
rect 1582 162 1592 164
rect 1582 158 1584 162
rect 1588 158 1592 162
rect 1582 156 1592 158
rect 1595 156 1607 164
rect 1610 162 1620 164
rect 1610 158 1614 162
rect 1618 158 1620 162
rect 1717 162 1719 166
rect 1723 162 1727 166
rect 1717 160 1727 162
rect 1730 160 1742 168
rect 1745 166 1755 168
rect 1745 162 1749 166
rect 1753 162 1755 166
rect 1745 160 1755 162
rect 1610 156 1620 158
rect 1649 118 1659 120
rect 1649 114 1651 118
rect 1655 114 1659 118
rect 1649 112 1659 114
rect 1662 112 1674 120
rect 1677 118 1687 120
rect 1677 114 1681 118
rect 1685 114 1687 118
rect 1677 112 1687 114
rect 1576 18 1586 20
rect 1576 14 1578 18
rect 1582 14 1586 18
rect 1576 12 1586 14
rect 1589 12 1601 20
rect 1604 18 1614 20
rect 1604 14 1608 18
rect 1612 14 1614 18
rect 1604 12 1614 14
rect 1618 18 1628 20
rect 1618 14 1620 18
rect 1624 14 1628 18
rect 1618 12 1628 14
rect 1630 18 1640 20
rect 1630 14 1634 18
rect 1638 14 1640 18
rect 1630 12 1640 14
rect 1863 199 1873 201
rect 1876 199 1888 207
rect 1891 205 1901 207
rect 1891 201 1895 205
rect 1899 201 1901 205
rect 1891 199 1901 201
rect 1931 170 1941 172
rect 1796 166 1806 168
rect 1796 162 1798 166
rect 1802 162 1806 166
rect 1796 160 1806 162
rect 1809 160 1821 168
rect 1824 166 1834 168
rect 1824 162 1828 166
rect 1832 162 1834 166
rect 1931 166 1933 170
rect 1937 166 1941 170
rect 1931 164 1941 166
rect 1944 164 1956 172
rect 1959 170 1969 172
rect 1959 166 1963 170
rect 1967 166 1969 170
rect 1959 164 1969 166
rect 1824 160 1834 162
rect 1863 122 1873 124
rect 1863 118 1865 122
rect 1869 118 1873 122
rect 1863 116 1873 118
rect 1876 116 1888 124
rect 1891 122 1901 124
rect 1891 118 1895 122
rect 1899 118 1901 122
rect 1891 116 1901 118
rect 1798 18 1808 20
rect 1798 14 1800 18
rect 1804 14 1808 18
rect 1798 12 1808 14
rect 1811 12 1823 20
rect 1826 18 1836 20
rect 1826 14 1830 18
rect 1834 14 1836 18
rect 1826 12 1836 14
rect 1840 18 1850 20
rect 1840 14 1842 18
rect 1846 14 1850 18
rect 1840 12 1850 14
rect 1852 18 1862 20
rect 1852 14 1856 18
rect 1860 14 1862 18
rect 1852 12 1862 14
rect 1910 18 1920 20
rect 1910 14 1912 18
rect 1916 14 1920 18
rect 1910 12 1920 14
rect 1923 18 1935 20
rect 1923 14 1926 18
rect 1930 14 1935 18
rect 1923 12 1935 14
rect 1938 18 1948 20
rect 1938 14 1942 18
rect 1946 14 1948 18
rect 1938 12 1948 14
rect 1952 18 1962 20
rect 1952 14 1954 18
rect 1958 14 1962 18
rect 1952 12 1962 14
rect 1964 18 1974 20
rect 1964 14 1968 18
rect 1972 14 1974 18
rect 1964 12 1974 14
<< pdiffusion >>
rect 307 246 317 248
rect 93 242 103 244
rect 93 238 95 242
rect 99 238 103 242
rect 93 236 103 238
rect 106 242 118 244
rect 106 238 110 242
rect 114 238 118 242
rect 106 236 118 238
rect 121 242 131 244
rect 121 238 125 242
rect 129 238 131 242
rect 307 242 309 246
rect 313 242 317 246
rect 307 240 317 242
rect 320 246 332 248
rect 320 242 324 246
rect 328 242 332 246
rect 320 240 332 242
rect 335 246 345 248
rect 335 242 339 246
rect 343 242 345 246
rect 814 245 824 247
rect 335 240 345 242
rect 600 241 610 243
rect 121 236 131 238
rect 600 237 602 241
rect 606 237 610 241
rect 600 235 610 237
rect 613 241 625 243
rect 613 237 617 241
rect 621 237 625 241
rect 613 235 625 237
rect 628 241 638 243
rect 628 237 632 241
rect 636 237 638 241
rect 814 241 816 245
rect 820 241 824 245
rect 814 239 824 241
rect 827 245 839 247
rect 827 241 831 245
rect 835 241 839 245
rect 827 239 839 241
rect 842 245 852 247
rect 842 241 846 245
rect 850 241 852 245
rect 1324 245 1334 247
rect 842 239 852 241
rect 1110 241 1120 243
rect 628 235 638 237
rect 26 203 36 205
rect 26 199 28 203
rect 32 199 36 203
rect 26 197 36 199
rect 39 203 51 205
rect 39 199 43 203
rect 47 199 51 203
rect 39 197 51 199
rect 54 203 64 205
rect 161 207 171 209
rect 54 199 58 203
rect 62 199 64 203
rect 54 197 64 199
rect 161 203 163 207
rect 167 203 171 207
rect 161 201 171 203
rect 174 207 186 209
rect 174 203 178 207
rect 182 203 186 207
rect 174 201 186 203
rect 189 207 199 209
rect 189 203 193 207
rect 197 203 199 207
rect 189 201 199 203
rect 240 207 250 209
rect 240 203 242 207
rect 246 203 250 207
rect 240 201 250 203
rect 253 207 265 209
rect 253 203 257 207
rect 261 203 265 207
rect 253 201 265 203
rect 268 207 278 209
rect 375 211 385 213
rect 268 203 272 207
rect 276 203 278 207
rect 268 201 278 203
rect 93 159 103 161
rect 93 155 95 159
rect 99 155 103 159
rect 93 153 103 155
rect 106 159 118 161
rect 106 155 110 159
rect 114 155 118 159
rect 106 153 118 155
rect 121 159 131 161
rect 121 155 125 159
rect 129 155 131 159
rect 121 153 131 155
rect 20 59 30 61
rect 20 55 22 59
rect 26 55 30 59
rect 20 53 30 55
rect 33 59 45 61
rect 33 55 37 59
rect 41 55 45 59
rect 33 53 45 55
rect 48 59 58 61
rect 48 55 52 59
rect 56 55 58 59
rect 48 53 58 55
rect 62 59 72 61
rect 62 55 64 59
rect 68 55 72 59
rect 62 53 72 55
rect 74 59 84 61
rect 74 55 78 59
rect 82 55 84 59
rect 74 53 84 55
rect 375 207 377 211
rect 381 207 385 211
rect 375 205 385 207
rect 388 211 400 213
rect 388 207 392 211
rect 396 207 400 211
rect 388 205 400 207
rect 403 211 413 213
rect 1110 237 1112 241
rect 1116 237 1120 241
rect 1110 235 1120 237
rect 1123 241 1135 243
rect 1123 237 1127 241
rect 1131 237 1135 241
rect 1123 235 1135 237
rect 1138 241 1148 243
rect 1138 237 1142 241
rect 1146 237 1148 241
rect 1324 241 1326 245
rect 1330 241 1334 245
rect 1324 239 1334 241
rect 1337 245 1349 247
rect 1337 241 1341 245
rect 1345 241 1349 245
rect 1337 239 1349 241
rect 1352 245 1362 247
rect 1352 241 1356 245
rect 1360 241 1362 245
rect 1863 245 1873 247
rect 1352 239 1362 241
rect 1649 241 1659 243
rect 1138 235 1148 237
rect 403 207 407 211
rect 411 207 413 211
rect 403 205 413 207
rect 533 202 543 204
rect 533 198 535 202
rect 539 198 543 202
rect 533 196 543 198
rect 546 202 558 204
rect 546 198 550 202
rect 554 198 558 202
rect 546 196 558 198
rect 561 202 571 204
rect 668 206 678 208
rect 561 198 565 202
rect 569 198 571 202
rect 561 196 571 198
rect 307 163 317 165
rect 307 159 309 163
rect 313 159 317 163
rect 307 157 317 159
rect 320 163 332 165
rect 320 159 324 163
rect 328 159 332 163
rect 320 157 332 159
rect 335 163 345 165
rect 335 159 339 163
rect 343 159 345 163
rect 335 157 345 159
rect 242 59 252 61
rect 242 55 244 59
rect 248 55 252 59
rect 242 53 252 55
rect 255 59 267 61
rect 255 55 259 59
rect 263 55 267 59
rect 255 53 267 55
rect 270 59 280 61
rect 270 55 274 59
rect 278 55 280 59
rect 270 53 280 55
rect 284 59 294 61
rect 284 55 286 59
rect 290 55 294 59
rect 284 53 294 55
rect 296 59 306 61
rect 296 55 300 59
rect 304 55 306 59
rect 296 53 306 55
rect 354 59 364 61
rect 354 55 356 59
rect 360 55 364 59
rect 354 53 364 55
rect 367 53 379 61
rect 382 59 392 61
rect 382 55 386 59
rect 390 55 392 59
rect 382 53 392 55
rect 396 59 406 61
rect 396 55 398 59
rect 402 55 406 59
rect 396 53 406 55
rect 408 59 418 61
rect 408 55 412 59
rect 416 55 418 59
rect 408 53 418 55
rect 668 202 670 206
rect 674 202 678 206
rect 668 200 678 202
rect 681 206 693 208
rect 681 202 685 206
rect 689 202 693 206
rect 681 200 693 202
rect 696 206 706 208
rect 696 202 700 206
rect 704 202 706 206
rect 696 200 706 202
rect 747 206 757 208
rect 747 202 749 206
rect 753 202 757 206
rect 747 200 757 202
rect 760 206 772 208
rect 760 202 764 206
rect 768 202 772 206
rect 760 200 772 202
rect 775 206 785 208
rect 1649 237 1651 241
rect 1655 237 1659 241
rect 1649 235 1659 237
rect 1662 241 1674 243
rect 1662 237 1666 241
rect 1670 237 1674 241
rect 1662 235 1674 237
rect 1677 241 1687 243
rect 1677 237 1681 241
rect 1685 237 1687 241
rect 1863 241 1865 245
rect 1869 241 1873 245
rect 1863 239 1873 241
rect 1876 245 1888 247
rect 1876 241 1880 245
rect 1884 241 1888 245
rect 1876 239 1888 241
rect 1891 245 1901 247
rect 1891 241 1895 245
rect 1899 241 1901 245
rect 1891 239 1901 241
rect 1677 235 1687 237
rect 882 210 892 212
rect 775 202 779 206
rect 783 202 785 206
rect 775 200 785 202
rect 600 158 610 160
rect 600 154 602 158
rect 606 154 610 158
rect 600 152 610 154
rect 613 158 625 160
rect 613 154 617 158
rect 621 154 625 158
rect 613 152 625 154
rect 628 158 638 160
rect 628 154 632 158
rect 636 154 638 158
rect 628 152 638 154
rect 527 58 537 60
rect 527 54 529 58
rect 533 54 537 58
rect 527 52 537 54
rect 540 58 552 60
rect 540 54 544 58
rect 548 54 552 58
rect 540 52 552 54
rect 555 58 565 60
rect 555 54 559 58
rect 563 54 565 58
rect 555 52 565 54
rect 569 58 579 60
rect 569 54 571 58
rect 575 54 579 58
rect 569 52 579 54
rect 581 58 591 60
rect 581 54 585 58
rect 589 54 591 58
rect 581 52 591 54
rect 882 206 884 210
rect 888 206 892 210
rect 882 204 892 206
rect 895 210 907 212
rect 895 206 899 210
rect 903 206 907 210
rect 895 204 907 206
rect 910 210 920 212
rect 910 206 914 210
rect 918 206 920 210
rect 910 204 920 206
rect 1043 202 1053 204
rect 1043 198 1045 202
rect 1049 198 1053 202
rect 1043 196 1053 198
rect 1056 202 1068 204
rect 1056 198 1060 202
rect 1064 198 1068 202
rect 1056 196 1068 198
rect 1071 202 1081 204
rect 1178 206 1188 208
rect 1071 198 1075 202
rect 1079 198 1081 202
rect 1071 196 1081 198
rect 814 162 824 164
rect 814 158 816 162
rect 820 158 824 162
rect 814 156 824 158
rect 827 162 839 164
rect 827 158 831 162
rect 835 158 839 162
rect 827 156 839 158
rect 842 162 852 164
rect 842 158 846 162
rect 850 158 852 162
rect 842 156 852 158
rect 749 58 759 60
rect 749 54 751 58
rect 755 54 759 58
rect 749 52 759 54
rect 762 58 774 60
rect 762 54 766 58
rect 770 54 774 58
rect 762 52 774 54
rect 777 58 787 60
rect 777 54 781 58
rect 785 54 787 58
rect 777 52 787 54
rect 791 58 801 60
rect 791 54 793 58
rect 797 54 801 58
rect 791 52 801 54
rect 803 58 813 60
rect 803 54 807 58
rect 811 54 813 58
rect 803 52 813 54
rect 861 58 871 60
rect 861 54 863 58
rect 867 54 871 58
rect 861 52 871 54
rect 874 52 886 60
rect 889 58 899 60
rect 889 54 893 58
rect 897 54 899 58
rect 889 52 899 54
rect 903 58 913 60
rect 903 54 905 58
rect 909 54 913 58
rect 903 52 913 54
rect 915 58 925 60
rect 915 54 919 58
rect 923 54 925 58
rect 915 52 925 54
rect 1178 202 1180 206
rect 1184 202 1188 206
rect 1178 200 1188 202
rect 1191 206 1203 208
rect 1191 202 1195 206
rect 1199 202 1203 206
rect 1191 200 1203 202
rect 1206 206 1216 208
rect 1206 202 1210 206
rect 1214 202 1216 206
rect 1206 200 1216 202
rect 1257 206 1267 208
rect 1257 202 1259 206
rect 1263 202 1267 206
rect 1257 200 1267 202
rect 1270 206 1282 208
rect 1270 202 1274 206
rect 1278 202 1282 206
rect 1270 200 1282 202
rect 1285 206 1295 208
rect 1392 210 1402 212
rect 1285 202 1289 206
rect 1293 202 1295 206
rect 1285 200 1295 202
rect 1110 158 1120 160
rect 1110 154 1112 158
rect 1116 154 1120 158
rect 1110 152 1120 154
rect 1123 158 1135 160
rect 1123 154 1127 158
rect 1131 154 1135 158
rect 1123 152 1135 154
rect 1138 158 1148 160
rect 1138 154 1142 158
rect 1146 154 1148 158
rect 1138 152 1148 154
rect 1037 58 1047 60
rect 1037 54 1039 58
rect 1043 54 1047 58
rect 1037 52 1047 54
rect 1050 58 1062 60
rect 1050 54 1054 58
rect 1058 54 1062 58
rect 1050 52 1062 54
rect 1065 58 1075 60
rect 1065 54 1069 58
rect 1073 54 1075 58
rect 1065 52 1075 54
rect 1079 58 1089 60
rect 1079 54 1081 58
rect 1085 54 1089 58
rect 1079 52 1089 54
rect 1091 58 1101 60
rect 1091 54 1095 58
rect 1099 54 1101 58
rect 1091 52 1101 54
rect 1392 206 1394 210
rect 1398 206 1402 210
rect 1392 204 1402 206
rect 1405 210 1417 212
rect 1405 206 1409 210
rect 1413 206 1417 210
rect 1405 204 1417 206
rect 1420 210 1430 212
rect 1420 206 1424 210
rect 1428 206 1430 210
rect 1420 204 1430 206
rect 1582 202 1592 204
rect 1582 198 1584 202
rect 1588 198 1592 202
rect 1582 196 1592 198
rect 1595 202 1607 204
rect 1595 198 1599 202
rect 1603 198 1607 202
rect 1595 196 1607 198
rect 1610 202 1620 204
rect 1717 206 1727 208
rect 1610 198 1614 202
rect 1618 198 1620 202
rect 1610 196 1620 198
rect 1324 162 1334 164
rect 1324 158 1326 162
rect 1330 158 1334 162
rect 1324 156 1334 158
rect 1337 162 1349 164
rect 1337 158 1341 162
rect 1345 158 1349 162
rect 1337 156 1349 158
rect 1352 162 1362 164
rect 1352 158 1356 162
rect 1360 158 1362 162
rect 1352 156 1362 158
rect 1259 58 1269 60
rect 1259 54 1261 58
rect 1265 54 1269 58
rect 1259 52 1269 54
rect 1272 58 1284 60
rect 1272 54 1276 58
rect 1280 54 1284 58
rect 1272 52 1284 54
rect 1287 58 1297 60
rect 1287 54 1291 58
rect 1295 54 1297 58
rect 1287 52 1297 54
rect 1301 58 1311 60
rect 1301 54 1303 58
rect 1307 54 1311 58
rect 1301 52 1311 54
rect 1313 58 1323 60
rect 1313 54 1317 58
rect 1321 54 1323 58
rect 1313 52 1323 54
rect 1371 58 1381 60
rect 1371 54 1373 58
rect 1377 54 1381 58
rect 1371 52 1381 54
rect 1384 52 1396 60
rect 1399 58 1409 60
rect 1399 54 1403 58
rect 1407 54 1409 58
rect 1399 52 1409 54
rect 1413 58 1423 60
rect 1413 54 1415 58
rect 1419 54 1423 58
rect 1413 52 1423 54
rect 1425 58 1435 60
rect 1425 54 1429 58
rect 1433 54 1435 58
rect 1425 52 1435 54
rect 1717 202 1719 206
rect 1723 202 1727 206
rect 1717 200 1727 202
rect 1730 206 1742 208
rect 1730 202 1734 206
rect 1738 202 1742 206
rect 1730 200 1742 202
rect 1745 206 1755 208
rect 1745 202 1749 206
rect 1753 202 1755 206
rect 1745 200 1755 202
rect 1796 206 1806 208
rect 1796 202 1798 206
rect 1802 202 1806 206
rect 1796 200 1806 202
rect 1809 206 1821 208
rect 1809 202 1813 206
rect 1817 202 1821 206
rect 1809 200 1821 202
rect 1824 206 1834 208
rect 1931 210 1941 212
rect 1824 202 1828 206
rect 1832 202 1834 206
rect 1824 200 1834 202
rect 1649 158 1659 160
rect 1649 154 1651 158
rect 1655 154 1659 158
rect 1649 152 1659 154
rect 1662 158 1674 160
rect 1662 154 1666 158
rect 1670 154 1674 158
rect 1662 152 1674 154
rect 1677 158 1687 160
rect 1677 154 1681 158
rect 1685 154 1687 158
rect 1677 152 1687 154
rect 1576 58 1586 60
rect 1576 54 1578 58
rect 1582 54 1586 58
rect 1576 52 1586 54
rect 1589 58 1601 60
rect 1589 54 1593 58
rect 1597 54 1601 58
rect 1589 52 1601 54
rect 1604 58 1614 60
rect 1604 54 1608 58
rect 1612 54 1614 58
rect 1604 52 1614 54
rect 1618 58 1628 60
rect 1618 54 1620 58
rect 1624 54 1628 58
rect 1618 52 1628 54
rect 1630 58 1640 60
rect 1630 54 1634 58
rect 1638 54 1640 58
rect 1630 52 1640 54
rect 1931 206 1933 210
rect 1937 206 1941 210
rect 1931 204 1941 206
rect 1944 210 1956 212
rect 1944 206 1948 210
rect 1952 206 1956 210
rect 1944 204 1956 206
rect 1959 210 1969 212
rect 1959 206 1963 210
rect 1967 206 1969 210
rect 1959 204 1969 206
rect 1863 162 1873 164
rect 1863 158 1865 162
rect 1869 158 1873 162
rect 1863 156 1873 158
rect 1876 162 1888 164
rect 1876 158 1880 162
rect 1884 158 1888 162
rect 1876 156 1888 158
rect 1891 162 1901 164
rect 1891 158 1895 162
rect 1899 158 1901 162
rect 1891 156 1901 158
rect 1798 58 1808 60
rect 1798 54 1800 58
rect 1804 54 1808 58
rect 1798 52 1808 54
rect 1811 58 1823 60
rect 1811 54 1815 58
rect 1819 54 1823 58
rect 1811 52 1823 54
rect 1826 58 1836 60
rect 1826 54 1830 58
rect 1834 54 1836 58
rect 1826 52 1836 54
rect 1840 58 1850 60
rect 1840 54 1842 58
rect 1846 54 1850 58
rect 1840 52 1850 54
rect 1852 58 1862 60
rect 1852 54 1856 58
rect 1860 54 1862 58
rect 1852 52 1862 54
rect 1910 58 1920 60
rect 1910 54 1912 58
rect 1916 54 1920 58
rect 1910 52 1920 54
rect 1923 52 1935 60
rect 1938 58 1948 60
rect 1938 54 1942 58
rect 1946 54 1948 58
rect 1938 52 1948 54
rect 1952 58 1962 60
rect 1952 54 1954 58
rect 1958 54 1962 58
rect 1952 52 1962 54
rect 1964 58 1974 60
rect 1964 54 1968 58
rect 1972 54 1974 58
rect 1964 52 1974 54
<< metal1 >>
rect -25 200 -21 301
rect -17 209 -13 301
rect 307 256 314 260
rect 318 256 333 260
rect 337 259 398 260
rect 337 256 397 259
rect 93 252 100 256
rect 104 252 119 256
rect 123 252 186 256
rect 95 242 99 252
rect 125 242 129 252
rect 110 229 114 238
rect 110 225 129 229
rect 16 221 91 225
rect 125 221 129 225
rect 180 221 184 252
rect 309 246 313 256
rect 339 246 343 256
rect 394 255 397 256
rect 324 233 328 242
rect 324 229 343 233
rect 230 225 305 229
rect 339 225 343 229
rect 394 225 398 255
rect -17 205 9 209
rect -25 196 -1 200
rect -36 186 -9 190
rect -13 99 -9 186
rect -5 174 -1 196
rect 5 182 9 205
rect 16 182 21 221
rect 87 217 113 221
rect 125 217 145 221
rect 161 217 168 221
rect 172 217 187 221
rect 191 217 201 221
rect 24 213 33 217
rect 37 213 52 217
rect 56 213 61 217
rect 28 203 32 213
rect 58 203 62 213
rect 78 209 98 213
rect 43 190 47 199
rect 43 186 62 190
rect 58 182 62 186
rect 78 182 82 209
rect 125 202 129 217
rect 95 190 99 198
rect 93 186 100 190
rect 104 186 121 190
rect 125 186 129 190
rect 141 186 145 217
rect 163 207 167 217
rect 193 207 197 217
rect 178 194 182 203
rect 178 190 197 194
rect 193 186 197 190
rect 230 186 235 225
rect 301 221 327 225
rect 339 221 359 225
rect 375 221 382 225
rect 386 221 401 225
rect 405 221 415 225
rect 238 217 247 221
rect 251 217 266 221
rect 270 217 275 221
rect 242 207 246 217
rect 272 207 276 217
rect 292 213 312 217
rect 257 194 261 203
rect 257 190 276 194
rect 272 186 276 190
rect 292 186 296 213
rect 339 206 343 221
rect 309 194 313 202
rect 307 190 314 194
rect 318 190 335 194
rect 339 190 343 194
rect 355 190 359 221
rect 377 211 381 221
rect 407 211 411 221
rect 392 198 396 207
rect 482 199 486 300
rect 490 208 494 300
rect 814 255 821 259
rect 825 255 840 259
rect 844 258 905 259
rect 844 255 904 258
rect 600 251 607 255
rect 611 251 626 255
rect 630 251 693 255
rect 602 241 606 251
rect 632 241 636 251
rect 617 228 621 237
rect 617 224 636 228
rect 523 220 598 224
rect 632 220 636 224
rect 687 220 691 251
rect 816 245 820 255
rect 846 245 850 255
rect 901 254 904 255
rect 831 232 835 241
rect 831 228 850 232
rect 737 224 812 228
rect 846 224 850 228
rect 901 224 905 254
rect 490 204 516 208
rect 392 194 411 198
rect 482 195 506 199
rect 407 190 411 194
rect 355 186 395 190
rect 407 186 440 190
rect 141 182 181 186
rect 193 184 260 186
rect 193 182 205 184
rect 5 181 46 182
rect 5 178 8 181
rect 12 178 46 181
rect 58 178 82 182
rect -5 172 31 174
rect -1 170 31 172
rect 18 143 23 170
rect 58 163 62 178
rect 28 151 32 159
rect 26 147 33 151
rect 37 147 54 151
rect 58 147 63 151
rect 18 139 73 143
rect 68 130 73 139
rect 78 138 82 178
rect 141 174 166 178
rect 94 169 100 173
rect 104 169 119 173
rect 123 169 131 173
rect 95 159 99 169
rect 125 159 129 169
rect 110 146 114 155
rect 110 142 129 146
rect 125 138 129 142
rect 141 138 145 174
rect 193 167 197 182
rect 209 182 260 184
rect 272 182 296 186
rect 217 174 245 178
rect 163 155 167 163
rect 163 151 168 155
rect 172 151 189 155
rect 193 151 197 155
rect 78 134 113 138
rect 125 134 145 138
rect 68 126 98 130
rect 125 119 129 134
rect 95 107 99 115
rect 95 103 100 107
rect 104 103 121 107
rect 125 103 129 107
rect 217 99 221 174
rect 232 147 237 174
rect 272 167 276 182
rect 242 155 246 163
rect 240 151 247 155
rect 251 151 268 155
rect 272 151 277 155
rect 232 143 287 147
rect 282 134 287 143
rect 292 142 296 182
rect 355 178 380 182
rect 308 173 314 177
rect 318 173 333 177
rect 337 173 345 177
rect 309 163 313 173
rect 339 163 343 173
rect 324 150 328 159
rect 324 146 343 150
rect 339 142 343 146
rect 355 142 359 178
rect 407 171 411 186
rect 464 185 498 189
rect 464 176 468 185
rect 435 172 468 176
rect 377 159 381 167
rect 377 155 382 159
rect 386 155 403 159
rect 407 155 411 159
rect 292 138 327 142
rect 339 138 359 142
rect 282 130 312 134
rect 339 123 343 138
rect 309 111 313 119
rect 309 107 314 111
rect 318 107 335 111
rect 339 107 343 111
rect -13 97 221 99
rect -13 95 217 97
rect 18 69 27 73
rect 31 69 46 73
rect 50 69 64 73
rect 68 69 78 73
rect 82 69 249 73
rect 253 69 268 73
rect 272 69 286 73
rect 290 69 300 73
rect 304 69 361 73
rect 365 69 380 73
rect 384 69 398 73
rect 402 69 412 73
rect 416 69 420 76
rect 22 59 26 69
rect 52 59 56 69
rect 64 59 68 69
rect 244 59 248 69
rect 274 59 278 69
rect 286 59 290 69
rect 356 59 360 69
rect 398 59 402 69
rect 37 46 41 55
rect 20 42 29 46
rect 37 42 56 46
rect 25 38 29 42
rect 52 38 56 42
rect 78 40 82 55
rect 259 46 263 55
rect 242 42 251 46
rect 259 42 278 46
rect 25 34 40 38
rect 52 34 68 38
rect 78 36 84 40
rect 247 38 251 42
rect 274 38 278 42
rect 300 40 304 55
rect 354 42 375 46
rect 20 26 25 30
rect 52 19 56 34
rect 78 19 82 36
rect 247 34 262 38
rect 274 34 290 38
rect 300 36 306 40
rect 386 38 390 55
rect 412 40 416 55
rect 435 40 439 172
rect 494 98 498 185
rect 502 173 506 195
rect 512 181 516 204
rect 523 181 528 220
rect 594 216 620 220
rect 632 216 652 220
rect 668 216 675 220
rect 679 216 694 220
rect 698 216 708 220
rect 531 212 540 216
rect 544 212 559 216
rect 563 212 568 216
rect 535 202 539 212
rect 565 202 569 212
rect 585 208 605 212
rect 550 189 554 198
rect 550 185 569 189
rect 565 181 569 185
rect 585 181 589 208
rect 632 201 636 216
rect 602 189 606 197
rect 600 185 607 189
rect 611 185 628 189
rect 632 185 636 189
rect 648 185 652 216
rect 670 206 674 216
rect 700 206 704 216
rect 685 193 689 202
rect 685 189 704 193
rect 700 185 704 189
rect 737 185 742 224
rect 808 220 834 224
rect 846 220 866 224
rect 882 220 889 224
rect 893 220 908 224
rect 912 220 922 224
rect 745 216 754 220
rect 758 216 773 220
rect 777 216 782 220
rect 749 206 753 216
rect 779 206 783 216
rect 799 212 819 216
rect 764 193 768 202
rect 764 189 783 193
rect 779 185 783 189
rect 799 185 803 212
rect 846 205 850 220
rect 816 193 820 201
rect 814 189 821 193
rect 825 189 842 193
rect 846 189 850 193
rect 862 189 866 220
rect 884 210 888 220
rect 914 210 918 220
rect 899 197 903 206
rect 992 199 996 300
rect 1000 208 1004 300
rect 1324 255 1331 259
rect 1335 255 1350 259
rect 1354 258 1415 259
rect 1354 255 1414 258
rect 1110 251 1117 255
rect 1121 251 1136 255
rect 1140 251 1203 255
rect 1112 241 1116 251
rect 1142 241 1146 251
rect 1127 228 1131 237
rect 1127 224 1146 228
rect 1033 220 1108 224
rect 1142 220 1146 224
rect 1197 220 1201 251
rect 1326 245 1330 255
rect 1356 245 1360 255
rect 1411 254 1414 255
rect 1341 232 1345 241
rect 1341 228 1360 232
rect 1247 224 1322 228
rect 1356 224 1360 228
rect 1411 224 1415 254
rect 1000 204 1026 208
rect 899 193 918 197
rect 992 195 1016 199
rect 914 189 918 193
rect 862 185 902 189
rect 914 185 947 189
rect 973 185 1008 189
rect 648 181 688 185
rect 700 183 767 185
rect 700 181 712 183
rect 512 180 553 181
rect 512 177 515 180
rect 519 177 553 180
rect 565 177 589 181
rect 502 171 538 173
rect 506 169 538 171
rect 525 142 530 169
rect 565 162 569 177
rect 535 150 539 158
rect 533 146 540 150
rect 544 146 561 150
rect 565 146 570 150
rect 525 138 580 142
rect 575 129 580 138
rect 585 137 589 177
rect 648 173 673 177
rect 601 168 607 172
rect 611 168 626 172
rect 630 168 638 172
rect 602 158 606 168
rect 632 158 636 168
rect 617 145 621 154
rect 617 141 636 145
rect 632 137 636 141
rect 648 137 652 173
rect 700 166 704 181
rect 716 181 767 183
rect 779 181 803 185
rect 724 173 752 177
rect 670 154 674 162
rect 670 150 675 154
rect 679 150 696 154
rect 700 150 704 154
rect 585 133 620 137
rect 632 133 652 137
rect 575 125 605 129
rect 632 118 636 133
rect 602 106 606 114
rect 602 102 607 106
rect 611 102 628 106
rect 632 102 636 106
rect 724 98 728 173
rect 739 146 744 173
rect 779 166 783 181
rect 749 154 753 162
rect 747 150 754 154
rect 758 150 775 154
rect 779 150 784 154
rect 739 142 794 146
rect 789 133 794 142
rect 799 141 803 181
rect 862 177 887 181
rect 815 172 821 176
rect 825 172 840 176
rect 844 172 852 176
rect 816 162 820 172
rect 846 162 850 172
rect 831 149 835 158
rect 831 145 850 149
rect 846 141 850 145
rect 862 141 866 177
rect 914 170 918 185
rect 973 175 977 185
rect 942 171 977 175
rect 884 158 888 166
rect 884 154 889 158
rect 893 154 910 158
rect 914 154 918 158
rect 799 137 834 141
rect 846 137 866 141
rect 789 129 819 133
rect 846 122 850 137
rect 816 110 820 118
rect 816 106 821 110
rect 825 106 842 110
rect 846 106 850 110
rect 494 96 728 98
rect 494 94 724 96
rect 525 68 534 72
rect 538 68 553 72
rect 557 68 571 72
rect 575 68 585 72
rect 589 68 756 72
rect 760 68 775 72
rect 779 68 793 72
rect 797 68 807 72
rect 811 68 868 72
rect 872 68 887 72
rect 891 68 905 72
rect 909 68 919 72
rect 923 68 927 75
rect 529 58 533 68
rect 559 58 563 68
rect 571 58 575 68
rect 751 58 755 68
rect 781 58 785 68
rect 793 58 797 68
rect 863 58 867 68
rect 905 58 909 68
rect 544 45 548 54
rect 527 41 536 45
rect 544 41 563 45
rect 241 26 247 30
rect 274 19 278 34
rect 300 19 304 36
rect 370 34 402 38
rect 412 36 439 40
rect 532 37 536 41
rect 559 37 563 41
rect 585 39 589 54
rect 766 45 770 54
rect 749 41 758 45
rect 766 41 785 45
rect 354 26 359 30
rect 370 19 374 34
rect 412 19 416 36
rect 532 33 547 37
rect 559 33 575 37
rect 585 35 591 39
rect 754 37 758 41
rect 781 37 785 41
rect 807 39 811 54
rect 861 41 882 45
rect 527 25 532 29
rect 22 7 26 15
rect 64 7 68 15
rect 20 3 27 7
rect 31 3 48 7
rect 52 3 64 7
rect 68 3 79 7
rect 83 5 145 7
rect 244 7 248 15
rect 286 7 290 15
rect 356 7 360 15
rect 386 7 390 15
rect 559 18 563 33
rect 585 18 589 35
rect 754 33 769 37
rect 781 33 797 37
rect 807 35 813 39
rect 893 37 897 54
rect 919 39 923 54
rect 942 39 946 171
rect 1004 98 1008 185
rect 1012 173 1016 195
rect 1022 181 1026 204
rect 1033 181 1038 220
rect 1104 216 1130 220
rect 1142 216 1162 220
rect 1178 216 1185 220
rect 1189 216 1204 220
rect 1208 216 1218 220
rect 1041 212 1050 216
rect 1054 212 1069 216
rect 1073 212 1078 216
rect 1045 202 1049 212
rect 1075 202 1079 212
rect 1095 208 1115 212
rect 1060 189 1064 198
rect 1060 185 1079 189
rect 1075 181 1079 185
rect 1095 181 1099 208
rect 1142 201 1146 216
rect 1112 189 1116 197
rect 1110 185 1117 189
rect 1121 185 1138 189
rect 1142 185 1146 189
rect 1158 185 1162 216
rect 1180 206 1184 216
rect 1210 206 1214 216
rect 1195 193 1199 202
rect 1195 189 1214 193
rect 1210 185 1214 189
rect 1247 185 1252 224
rect 1318 220 1344 224
rect 1356 220 1376 224
rect 1392 220 1399 224
rect 1403 220 1418 224
rect 1422 220 1432 224
rect 1255 216 1264 220
rect 1268 216 1283 220
rect 1287 216 1292 220
rect 1259 206 1263 216
rect 1289 206 1293 216
rect 1309 212 1329 216
rect 1274 193 1278 202
rect 1274 189 1293 193
rect 1289 185 1293 189
rect 1309 185 1313 212
rect 1356 205 1360 220
rect 1326 193 1330 201
rect 1324 189 1331 193
rect 1335 189 1352 193
rect 1356 189 1360 193
rect 1372 189 1376 220
rect 1394 210 1398 220
rect 1424 210 1428 220
rect 1409 197 1413 206
rect 1531 199 1535 300
rect 1539 208 1543 300
rect 1863 255 1870 259
rect 1874 255 1889 259
rect 1893 258 1954 259
rect 1893 255 1953 258
rect 1649 251 1656 255
rect 1660 251 1675 255
rect 1679 251 1742 255
rect 1651 241 1655 251
rect 1681 241 1685 251
rect 1666 228 1670 237
rect 1666 224 1685 228
rect 1572 220 1647 224
rect 1681 220 1685 224
rect 1736 220 1740 251
rect 1865 245 1869 255
rect 1895 245 1899 255
rect 1950 254 1953 255
rect 1880 232 1884 241
rect 1880 228 1899 232
rect 1786 224 1861 228
rect 1895 224 1899 228
rect 1950 224 1954 254
rect 1539 204 1565 208
rect 1409 193 1428 197
rect 1531 195 1555 199
rect 1424 189 1428 193
rect 1372 185 1412 189
rect 1424 185 1457 189
rect 1511 185 1547 189
rect 1158 181 1198 185
rect 1210 183 1277 185
rect 1210 181 1222 183
rect 1022 180 1063 181
rect 1022 177 1025 180
rect 1029 177 1063 180
rect 1075 177 1099 181
rect 1012 171 1048 173
rect 1016 169 1048 171
rect 1035 142 1040 169
rect 1075 162 1079 177
rect 1045 150 1049 158
rect 1043 146 1050 150
rect 1054 146 1071 150
rect 1075 146 1080 150
rect 1035 138 1090 142
rect 1085 129 1090 138
rect 1095 137 1099 177
rect 1158 173 1183 177
rect 1111 168 1117 172
rect 1121 168 1136 172
rect 1140 168 1148 172
rect 1112 158 1116 168
rect 1142 158 1146 168
rect 1127 145 1131 154
rect 1127 141 1146 145
rect 1142 137 1146 141
rect 1158 137 1162 173
rect 1210 166 1214 181
rect 1226 181 1277 183
rect 1289 181 1313 185
rect 1234 173 1262 177
rect 1180 154 1184 162
rect 1180 150 1185 154
rect 1189 150 1206 154
rect 1210 150 1214 154
rect 1095 133 1130 137
rect 1142 133 1162 137
rect 1085 125 1115 129
rect 1142 118 1146 133
rect 1112 106 1116 114
rect 1112 102 1117 106
rect 1121 102 1138 106
rect 1142 102 1146 106
rect 1234 98 1238 173
rect 1249 146 1254 173
rect 1289 166 1293 181
rect 1259 154 1263 162
rect 1257 150 1264 154
rect 1268 150 1285 154
rect 1289 150 1294 154
rect 1249 142 1304 146
rect 1299 133 1304 142
rect 1309 141 1313 181
rect 1372 177 1397 181
rect 1325 172 1331 176
rect 1335 172 1350 176
rect 1354 172 1362 176
rect 1326 162 1330 172
rect 1356 162 1360 172
rect 1341 149 1345 158
rect 1341 145 1360 149
rect 1356 141 1360 145
rect 1372 141 1376 177
rect 1424 170 1428 185
rect 1511 175 1515 185
rect 1452 171 1515 175
rect 1394 158 1398 166
rect 1394 154 1399 158
rect 1403 154 1420 158
rect 1424 154 1428 158
rect 1309 137 1344 141
rect 1356 137 1376 141
rect 1299 129 1329 133
rect 1356 122 1360 137
rect 1326 110 1330 118
rect 1326 106 1331 110
rect 1335 106 1352 110
rect 1356 106 1360 110
rect 1004 96 1238 98
rect 1004 94 1234 96
rect 1035 68 1044 72
rect 1048 68 1063 72
rect 1067 68 1081 72
rect 1085 68 1095 72
rect 1099 68 1266 72
rect 1270 68 1285 72
rect 1289 68 1303 72
rect 1307 68 1317 72
rect 1321 68 1378 72
rect 1382 68 1397 72
rect 1401 68 1415 72
rect 1419 68 1429 72
rect 1433 68 1437 75
rect 1039 58 1043 68
rect 1069 58 1073 68
rect 1081 58 1085 68
rect 1261 58 1265 68
rect 1291 58 1295 68
rect 1303 58 1307 68
rect 1373 58 1377 68
rect 1415 58 1419 68
rect 1054 45 1058 54
rect 1037 41 1046 45
rect 1054 41 1073 45
rect 748 25 754 29
rect 781 18 785 33
rect 807 18 811 35
rect 877 33 909 37
rect 919 35 946 39
rect 1042 37 1046 41
rect 1069 37 1073 41
rect 1095 39 1099 54
rect 1276 45 1280 54
rect 1259 41 1268 45
rect 1276 41 1295 45
rect 861 25 866 29
rect 877 18 881 33
rect 919 18 923 35
rect 1042 33 1057 37
rect 1069 33 1085 37
rect 1095 35 1101 39
rect 1264 37 1268 41
rect 1291 37 1295 41
rect 1317 39 1321 54
rect 1371 41 1392 45
rect 1037 25 1042 29
rect 1069 18 1073 33
rect 1095 18 1099 35
rect 1264 33 1279 37
rect 1291 33 1307 37
rect 1317 35 1323 39
rect 1403 37 1407 54
rect 1429 39 1433 54
rect 1452 39 1456 171
rect 1543 98 1547 185
rect 1551 173 1555 195
rect 1561 181 1565 204
rect 1572 181 1577 220
rect 1643 216 1669 220
rect 1681 216 1701 220
rect 1717 216 1724 220
rect 1728 216 1743 220
rect 1747 216 1757 220
rect 1580 212 1589 216
rect 1593 212 1608 216
rect 1612 212 1617 216
rect 1584 202 1588 212
rect 1614 202 1618 212
rect 1634 208 1654 212
rect 1599 189 1603 198
rect 1599 185 1618 189
rect 1614 181 1618 185
rect 1634 181 1638 208
rect 1681 201 1685 216
rect 1651 189 1655 197
rect 1649 185 1656 189
rect 1660 185 1677 189
rect 1681 185 1685 189
rect 1697 185 1701 216
rect 1719 206 1723 216
rect 1749 206 1753 216
rect 1734 193 1738 202
rect 1734 189 1753 193
rect 1749 185 1753 189
rect 1786 185 1791 224
rect 1857 220 1883 224
rect 1895 220 1915 224
rect 1931 220 1938 224
rect 1942 220 1957 224
rect 1961 220 1971 224
rect 1794 216 1803 220
rect 1807 216 1822 220
rect 1826 216 1831 220
rect 1798 206 1802 216
rect 1828 206 1832 216
rect 1848 212 1868 216
rect 1813 193 1817 202
rect 1813 189 1832 193
rect 1828 185 1832 189
rect 1848 185 1852 212
rect 1895 205 1899 220
rect 1865 193 1869 201
rect 1863 189 1870 193
rect 1874 189 1891 193
rect 1895 189 1899 193
rect 1911 189 1915 220
rect 1933 210 1937 220
rect 1963 210 1967 220
rect 1948 197 1952 206
rect 1948 193 1967 197
rect 1963 189 1967 193
rect 1911 185 1951 189
rect 1963 185 1996 189
rect 1697 181 1737 185
rect 1749 183 1816 185
rect 1749 181 1761 183
rect 1561 180 1602 181
rect 1561 177 1564 180
rect 1568 177 1602 180
rect 1614 177 1638 181
rect 1551 171 1587 173
rect 1555 169 1587 171
rect 1574 142 1579 169
rect 1614 162 1618 177
rect 1584 150 1588 158
rect 1582 146 1589 150
rect 1593 146 1610 150
rect 1614 146 1619 150
rect 1574 138 1629 142
rect 1624 129 1629 138
rect 1634 137 1638 177
rect 1697 173 1722 177
rect 1650 168 1656 172
rect 1660 168 1675 172
rect 1679 168 1687 172
rect 1651 158 1655 168
rect 1681 158 1685 168
rect 1666 145 1670 154
rect 1666 141 1685 145
rect 1681 137 1685 141
rect 1697 137 1701 173
rect 1749 166 1753 181
rect 1765 181 1816 183
rect 1828 181 1852 185
rect 1773 173 1801 177
rect 1719 154 1723 162
rect 1719 150 1724 154
rect 1728 150 1745 154
rect 1749 150 1753 154
rect 1634 133 1669 137
rect 1681 133 1701 137
rect 1624 125 1654 129
rect 1681 118 1685 133
rect 1651 106 1655 114
rect 1651 102 1656 106
rect 1660 102 1677 106
rect 1681 102 1685 106
rect 1773 98 1777 173
rect 1788 146 1793 173
rect 1828 166 1832 181
rect 1798 154 1802 162
rect 1796 150 1803 154
rect 1807 150 1824 154
rect 1828 150 1833 154
rect 1788 142 1843 146
rect 1838 133 1843 142
rect 1848 141 1852 181
rect 1911 177 1936 181
rect 1864 172 1870 176
rect 1874 172 1889 176
rect 1893 172 1901 176
rect 1865 162 1869 172
rect 1895 162 1899 172
rect 1880 149 1884 158
rect 1880 145 1899 149
rect 1895 141 1899 145
rect 1911 141 1915 177
rect 1963 170 1967 185
rect 1991 171 1998 175
rect 1933 158 1937 166
rect 1933 154 1938 158
rect 1942 154 1959 158
rect 1963 154 1967 158
rect 1848 137 1883 141
rect 1895 137 1915 141
rect 1838 129 1868 133
rect 1895 122 1899 137
rect 1865 110 1869 118
rect 1865 106 1870 110
rect 1874 106 1891 110
rect 1895 106 1899 110
rect 1543 96 1777 98
rect 1543 94 1773 96
rect 1574 68 1583 72
rect 1587 68 1602 72
rect 1606 68 1620 72
rect 1624 68 1634 72
rect 1638 68 1805 72
rect 1809 68 1824 72
rect 1828 68 1842 72
rect 1846 68 1856 72
rect 1860 68 1917 72
rect 1921 68 1936 72
rect 1940 68 1954 72
rect 1958 68 1968 72
rect 1972 68 1976 75
rect 1578 58 1582 68
rect 1608 58 1612 68
rect 1620 58 1624 68
rect 1800 58 1804 68
rect 1830 58 1834 68
rect 1842 58 1846 68
rect 1912 58 1916 68
rect 1954 58 1958 68
rect 1593 45 1597 54
rect 1576 41 1585 45
rect 1593 41 1612 45
rect 1258 25 1264 29
rect 1291 18 1295 33
rect 1317 18 1321 35
rect 1387 33 1419 37
rect 1429 35 1456 39
rect 1581 37 1585 41
rect 1608 37 1612 41
rect 1634 39 1638 54
rect 1815 45 1819 54
rect 1798 41 1807 45
rect 1815 41 1834 45
rect 1371 25 1376 29
rect 1387 18 1391 33
rect 1429 18 1433 35
rect 1581 33 1596 37
rect 1608 33 1624 37
rect 1634 35 1640 39
rect 1803 37 1807 41
rect 1830 37 1834 41
rect 1856 39 1860 54
rect 1910 41 1931 45
rect 1576 25 1581 29
rect 1608 18 1612 33
rect 1634 18 1638 35
rect 1803 33 1818 37
rect 1830 33 1846 37
rect 1856 35 1862 39
rect 1942 37 1946 54
rect 1968 39 1972 54
rect 1991 39 1995 171
rect 1797 25 1803 29
rect 1830 18 1834 33
rect 1856 18 1860 35
rect 1926 33 1958 37
rect 1968 35 1995 39
rect 1912 25 1915 29
rect 1926 18 1930 33
rect 1968 18 1972 35
rect 398 7 402 15
rect 149 5 249 7
rect 83 3 249 5
rect 253 3 270 7
rect 274 3 286 7
rect 290 3 301 7
rect 305 3 361 7
rect 365 3 382 7
rect 386 3 398 7
rect 402 3 413 7
rect 417 3 422 7
rect 523 6 524 7
rect 529 6 533 14
rect 571 6 575 14
rect 523 2 534 6
rect 538 2 555 6
rect 559 2 571 6
rect 575 2 586 6
rect 590 4 652 6
rect 751 6 755 14
rect 793 6 797 14
rect 863 6 867 14
rect 893 6 897 14
rect 905 6 909 14
rect 1039 6 1043 14
rect 1081 6 1085 14
rect 656 4 756 6
rect 590 2 756 4
rect 760 2 777 6
rect 781 2 793 6
rect 797 2 808 6
rect 812 2 868 6
rect 872 2 889 6
rect 893 2 905 6
rect 909 2 920 6
rect 924 2 925 6
rect 1039 2 1044 6
rect 1048 2 1065 6
rect 1069 2 1081 6
rect 1085 2 1096 6
rect 1100 4 1162 6
rect 1261 6 1265 14
rect 1303 6 1307 14
rect 1373 6 1377 14
rect 1403 6 1407 14
rect 1415 6 1419 14
rect 1578 6 1582 14
rect 1620 6 1624 14
rect 1166 4 1266 6
rect 1100 2 1266 4
rect 1270 2 1287 6
rect 1291 2 1303 6
rect 1307 2 1318 6
rect 1322 2 1378 6
rect 1382 2 1399 6
rect 1403 2 1415 6
rect 1419 2 1430 6
rect 1434 2 1435 6
rect 1578 2 1583 6
rect 1587 2 1604 6
rect 1608 2 1620 6
rect 1624 2 1635 6
rect 1639 4 1701 6
rect 1800 6 1804 14
rect 1842 6 1846 14
rect 1912 6 1916 14
rect 1942 6 1946 14
rect 1954 6 1958 14
rect 1705 4 1805 6
rect 1639 2 1805 4
rect 1809 2 1826 6
rect 1830 2 1842 6
rect 1846 2 1857 6
rect 1861 2 1917 6
rect 1921 2 1938 6
rect 1942 2 1954 6
rect 1958 2 1969 6
rect 1973 2 1976 6
<< metal2 >>
rect 277 256 303 260
rect 63 252 89 256
rect 190 252 281 256
rect 401 255 426 259
rect 784 255 810 259
rect 63 217 67 252
rect 277 221 281 252
rect 422 251 426 255
rect 570 251 596 255
rect 697 251 788 255
rect 908 254 933 258
rect 1294 255 1320 259
rect 422 247 574 251
rect 279 217 289 221
rect 65 213 75 217
rect 71 173 75 213
rect 71 169 90 173
rect 67 147 77 151
rect 73 107 77 147
rect 133 107 137 190
rect 285 177 289 217
rect 285 173 304 177
rect 157 151 159 155
rect 281 151 291 155
rect 157 107 161 151
rect 287 118 291 151
rect 257 114 291 118
rect 257 107 261 114
rect 287 111 291 114
rect 347 111 351 194
rect 371 155 373 159
rect 422 156 426 247
rect 570 216 574 247
rect 784 220 788 251
rect 929 246 933 254
rect 1080 251 1106 255
rect 1207 251 1298 255
rect 1418 254 1443 258
rect 1833 255 1859 259
rect 1080 246 1084 251
rect 929 242 1084 246
rect 786 216 796 220
rect 572 212 582 216
rect 578 172 582 212
rect 578 168 597 172
rect 371 111 375 155
rect 287 107 305 111
rect 347 107 375 111
rect 416 152 426 156
rect 73 103 91 107
rect 133 103 261 107
rect 145 9 149 103
rect 416 80 420 152
rect 574 146 584 150
rect 580 106 584 146
rect 640 106 644 189
rect 792 176 796 216
rect 792 172 811 176
rect 664 150 666 154
rect 788 150 798 154
rect 664 106 668 150
rect 794 117 798 150
rect 764 113 798 117
rect 764 106 768 113
rect 794 110 798 113
rect 854 110 858 193
rect 878 154 880 158
rect 929 155 933 242
rect 1080 216 1084 242
rect 1294 220 1298 251
rect 1439 243 1443 254
rect 1619 251 1645 255
rect 1746 251 1837 255
rect 1957 254 1982 258
rect 1619 243 1623 251
rect 1439 239 1624 243
rect 1296 216 1306 220
rect 1082 212 1092 216
rect 1088 172 1092 212
rect 1088 168 1107 172
rect 878 110 882 154
rect 794 106 812 110
rect 854 106 882 110
rect 923 151 933 155
rect 580 102 598 106
rect 640 102 768 106
rect 652 8 656 102
rect 923 79 927 151
rect 1084 146 1094 150
rect 1090 106 1094 146
rect 1150 106 1154 189
rect 1302 176 1306 216
rect 1302 172 1321 176
rect 1174 150 1176 154
rect 1298 150 1308 154
rect 1174 106 1178 150
rect 1304 117 1308 150
rect 1274 113 1308 117
rect 1274 106 1278 113
rect 1304 110 1308 113
rect 1364 110 1368 193
rect 1388 154 1390 158
rect 1439 155 1443 239
rect 1619 216 1623 239
rect 1833 220 1837 251
rect 1835 216 1845 220
rect 1621 212 1631 216
rect 1627 172 1631 212
rect 1627 168 1646 172
rect 1388 110 1392 154
rect 1304 106 1322 110
rect 1364 106 1392 110
rect 1433 151 1443 155
rect 1090 102 1108 106
rect 1150 102 1278 106
rect 426 3 519 7
rect 517 2 519 3
rect 1162 8 1166 102
rect 1433 79 1437 151
rect 1623 146 1633 150
rect 1629 106 1633 146
rect 1689 106 1693 189
rect 1841 176 1845 216
rect 1841 172 1860 176
rect 1713 150 1715 154
rect 1837 150 1847 154
rect 1713 106 1717 150
rect 1843 117 1847 150
rect 1813 113 1847 117
rect 1813 106 1817 113
rect 1843 110 1847 113
rect 1903 110 1907 193
rect 1927 154 1929 158
rect 1978 155 1982 254
rect 1927 110 1931 154
rect 1843 106 1861 110
rect 1903 106 1931 110
rect 1972 151 1982 155
rect 1629 102 1647 106
rect 1689 102 1817 106
rect 929 2 1035 6
rect 1701 8 1705 102
rect 1972 79 1976 151
rect 1439 2 1574 6
<< ntransistor >>
rect 103 196 106 204
rect 118 196 121 204
rect 36 157 39 165
rect 51 157 54 165
rect 171 161 174 169
rect 186 161 189 169
rect 103 113 106 121
rect 118 113 121 121
rect 30 13 33 21
rect 45 13 48 21
rect 72 13 74 21
rect 317 200 320 208
rect 332 200 335 208
rect 250 161 253 169
rect 265 161 268 169
rect 385 165 388 173
rect 400 165 403 173
rect 317 117 320 125
rect 332 117 335 125
rect 252 13 255 21
rect 267 13 270 21
rect 294 13 296 21
rect 364 13 367 21
rect 379 13 382 21
rect 406 13 408 21
rect 610 195 613 203
rect 625 195 628 203
rect 543 156 546 164
rect 558 156 561 164
rect 678 160 681 168
rect 693 160 696 168
rect 610 112 613 120
rect 625 112 628 120
rect 537 12 540 20
rect 552 12 555 20
rect 579 12 581 20
rect 824 199 827 207
rect 839 199 842 207
rect 757 160 760 168
rect 772 160 775 168
rect 892 164 895 172
rect 907 164 910 172
rect 824 116 827 124
rect 839 116 842 124
rect 759 12 762 20
rect 774 12 777 20
rect 801 12 803 20
rect 871 12 874 20
rect 886 12 889 20
rect 913 12 915 20
rect 1120 195 1123 203
rect 1135 195 1138 203
rect 1053 156 1056 164
rect 1068 156 1071 164
rect 1188 160 1191 168
rect 1203 160 1206 168
rect 1120 112 1123 120
rect 1135 112 1138 120
rect 1047 12 1050 20
rect 1062 12 1065 20
rect 1089 12 1091 20
rect 1334 199 1337 207
rect 1349 199 1352 207
rect 1267 160 1270 168
rect 1282 160 1285 168
rect 1402 164 1405 172
rect 1417 164 1420 172
rect 1334 116 1337 124
rect 1349 116 1352 124
rect 1269 12 1272 20
rect 1284 12 1287 20
rect 1311 12 1313 20
rect 1381 12 1384 20
rect 1396 12 1399 20
rect 1423 12 1425 20
rect 1659 195 1662 203
rect 1674 195 1677 203
rect 1592 156 1595 164
rect 1607 156 1610 164
rect 1727 160 1730 168
rect 1742 160 1745 168
rect 1659 112 1662 120
rect 1674 112 1677 120
rect 1586 12 1589 20
rect 1601 12 1604 20
rect 1628 12 1630 20
rect 1873 199 1876 207
rect 1888 199 1891 207
rect 1806 160 1809 168
rect 1821 160 1824 168
rect 1941 164 1944 172
rect 1956 164 1959 172
rect 1873 116 1876 124
rect 1888 116 1891 124
rect 1808 12 1811 20
rect 1823 12 1826 20
rect 1850 12 1852 20
rect 1920 12 1923 20
rect 1935 12 1938 20
rect 1962 12 1964 20
<< ptransistor >>
rect 103 236 106 244
rect 118 236 121 244
rect 317 240 320 248
rect 332 240 335 248
rect 610 235 613 243
rect 625 235 628 243
rect 824 239 827 247
rect 839 239 842 247
rect 36 197 39 205
rect 51 197 54 205
rect 171 201 174 209
rect 186 201 189 209
rect 250 201 253 209
rect 265 201 268 209
rect 103 153 106 161
rect 118 153 121 161
rect 30 53 33 61
rect 45 53 48 61
rect 72 53 74 61
rect 385 205 388 213
rect 400 205 403 213
rect 1120 235 1123 243
rect 1135 235 1138 243
rect 1334 239 1337 247
rect 1349 239 1352 247
rect 543 196 546 204
rect 558 196 561 204
rect 317 157 320 165
rect 332 157 335 165
rect 252 53 255 61
rect 267 53 270 61
rect 294 53 296 61
rect 364 53 367 61
rect 379 53 382 61
rect 406 53 408 61
rect 678 200 681 208
rect 693 200 696 208
rect 757 200 760 208
rect 772 200 775 208
rect 1659 235 1662 243
rect 1674 235 1677 243
rect 1873 239 1876 247
rect 1888 239 1891 247
rect 610 152 613 160
rect 625 152 628 160
rect 537 52 540 60
rect 552 52 555 60
rect 579 52 581 60
rect 892 204 895 212
rect 907 204 910 212
rect 1053 196 1056 204
rect 1068 196 1071 204
rect 824 156 827 164
rect 839 156 842 164
rect 759 52 762 60
rect 774 52 777 60
rect 801 52 803 60
rect 871 52 874 60
rect 886 52 889 60
rect 913 52 915 60
rect 1188 200 1191 208
rect 1203 200 1206 208
rect 1267 200 1270 208
rect 1282 200 1285 208
rect 1120 152 1123 160
rect 1135 152 1138 160
rect 1047 52 1050 60
rect 1062 52 1065 60
rect 1089 52 1091 60
rect 1402 204 1405 212
rect 1417 204 1420 212
rect 1592 196 1595 204
rect 1607 196 1610 204
rect 1334 156 1337 164
rect 1349 156 1352 164
rect 1269 52 1272 60
rect 1284 52 1287 60
rect 1311 52 1313 60
rect 1381 52 1384 60
rect 1396 52 1399 60
rect 1423 52 1425 60
rect 1727 200 1730 208
rect 1742 200 1745 208
rect 1806 200 1809 208
rect 1821 200 1824 208
rect 1659 152 1662 160
rect 1674 152 1677 160
rect 1586 52 1589 60
rect 1601 52 1604 60
rect 1628 52 1630 60
rect 1941 204 1944 212
rect 1956 204 1959 212
rect 1873 156 1876 164
rect 1888 156 1891 164
rect 1808 52 1811 60
rect 1823 52 1826 60
rect 1850 52 1852 60
rect 1920 52 1923 60
rect 1935 52 1938 60
rect 1962 52 1964 60
<< polycontact >>
rect 113 217 117 221
rect 327 221 331 225
rect 98 209 102 213
rect 312 213 316 217
rect 8 177 12 181
rect -5 168 -1 172
rect 46 178 50 182
rect 181 182 185 186
rect 31 170 35 174
rect 166 174 170 178
rect 205 180 209 184
rect 113 134 117 138
rect 98 126 102 130
rect 16 42 20 46
rect 40 34 44 38
rect 68 34 72 38
rect 16 26 20 30
rect 25 26 29 30
rect 84 36 88 40
rect 620 216 624 220
rect 834 220 838 224
rect 605 208 609 212
rect 260 182 264 186
rect 819 212 823 216
rect 395 186 399 190
rect 440 186 444 190
rect 245 174 249 178
rect 380 178 384 182
rect 327 138 331 142
rect 312 130 316 134
rect 217 93 221 97
rect 238 42 242 46
rect 262 34 266 38
rect 290 34 294 38
rect 237 26 241 30
rect 247 26 251 30
rect 350 42 354 46
rect 306 36 311 40
rect 375 42 379 46
rect 350 26 354 30
rect 359 26 363 30
rect 402 34 406 38
rect 515 176 519 180
rect 502 167 506 171
rect 1130 216 1134 220
rect 1344 220 1348 224
rect 553 177 557 181
rect 688 181 692 185
rect 538 169 542 173
rect 673 173 677 177
rect 712 179 716 183
rect 620 133 624 137
rect 605 125 609 129
rect 523 41 527 45
rect 547 33 551 37
rect 575 33 579 37
rect 523 25 527 29
rect 532 25 536 29
rect 591 35 595 39
rect 1115 208 1119 212
rect 767 181 771 185
rect 1329 212 1333 216
rect 902 185 906 189
rect 947 185 951 189
rect 752 173 756 177
rect 887 177 891 181
rect 834 137 838 141
rect 819 129 823 133
rect 724 92 728 96
rect 745 41 749 45
rect 769 33 773 37
rect 797 33 801 37
rect 744 25 748 29
rect 754 25 758 29
rect 857 41 861 45
rect 813 35 818 39
rect 882 41 886 45
rect 857 25 861 29
rect 866 25 870 29
rect 909 33 913 37
rect 1025 176 1029 180
rect 1012 167 1016 171
rect 1669 216 1673 220
rect 1883 220 1887 224
rect 1063 177 1067 181
rect 1198 181 1202 185
rect 1048 169 1052 173
rect 1183 173 1187 177
rect 1222 179 1226 183
rect 1130 133 1134 137
rect 1115 125 1119 129
rect 1033 41 1037 45
rect 1057 33 1061 37
rect 1085 33 1089 37
rect 1033 25 1037 29
rect 1042 25 1046 29
rect 1101 35 1105 39
rect 1654 208 1658 212
rect 1277 181 1281 185
rect 1868 212 1872 216
rect 1412 185 1416 189
rect 1457 185 1461 189
rect 1262 173 1266 177
rect 1397 177 1401 181
rect 1344 137 1348 141
rect 1329 129 1333 133
rect 1234 92 1238 96
rect 1255 41 1259 45
rect 1279 33 1283 37
rect 1307 33 1311 37
rect 1254 25 1258 29
rect 1264 25 1268 29
rect 1367 41 1371 45
rect 1323 35 1328 39
rect 1392 41 1396 45
rect 1367 25 1371 29
rect 1376 25 1380 29
rect 1419 33 1423 37
rect 1564 176 1568 180
rect 1551 167 1555 171
rect 1602 177 1606 181
rect 1737 181 1741 185
rect 1587 169 1591 173
rect 1722 173 1726 177
rect 1761 179 1765 183
rect 1669 133 1673 137
rect 1654 125 1658 129
rect 1572 41 1576 45
rect 1596 33 1600 37
rect 1624 33 1628 37
rect 1572 25 1576 29
rect 1581 25 1585 29
rect 1640 35 1644 39
rect 1816 181 1820 185
rect 1951 185 1955 189
rect 1996 185 2000 189
rect 1801 173 1805 177
rect 1936 177 1940 181
rect 1998 171 2002 175
rect 1883 137 1887 141
rect 1868 129 1872 133
rect 1773 92 1777 96
rect 1794 41 1798 45
rect 1818 33 1822 37
rect 1846 33 1850 37
rect 1793 25 1797 29
rect 1803 25 1807 29
rect 1906 41 1910 45
rect 1862 35 1867 39
rect 1931 41 1935 45
rect 1908 25 1912 29
rect 1915 25 1919 29
rect 1958 33 1962 37
<< ndcontact >>
rect 95 198 99 202
rect 125 198 129 202
rect 309 202 313 206
rect 28 159 32 163
rect 58 159 62 163
rect 163 163 167 167
rect 193 163 197 167
rect 95 115 99 119
rect 125 115 129 119
rect 22 15 26 19
rect 52 15 56 19
rect 64 15 68 19
rect 78 15 82 19
rect 339 202 343 206
rect 602 197 606 201
rect 242 163 246 167
rect 272 163 276 167
rect 377 167 381 171
rect 407 167 411 171
rect 309 119 313 123
rect 339 119 343 123
rect 244 15 248 19
rect 274 15 278 19
rect 286 15 290 19
rect 300 15 304 19
rect 356 15 360 19
rect 370 15 374 19
rect 386 15 390 19
rect 398 15 402 19
rect 412 15 416 19
rect 632 197 636 201
rect 816 201 820 205
rect 535 158 539 162
rect 565 158 569 162
rect 670 162 674 166
rect 700 162 704 166
rect 602 114 606 118
rect 632 114 636 118
rect 529 14 533 18
rect 559 14 563 18
rect 571 14 575 18
rect 585 14 589 18
rect 846 201 850 205
rect 1112 197 1116 201
rect 749 162 753 166
rect 779 162 783 166
rect 884 166 888 170
rect 914 166 918 170
rect 816 118 820 122
rect 846 118 850 122
rect 751 14 755 18
rect 781 14 785 18
rect 793 14 797 18
rect 807 14 811 18
rect 863 14 867 18
rect 877 14 881 18
rect 893 14 897 18
rect 905 14 909 18
rect 919 14 923 18
rect 1142 197 1146 201
rect 1326 201 1330 205
rect 1045 158 1049 162
rect 1075 158 1079 162
rect 1180 162 1184 166
rect 1210 162 1214 166
rect 1112 114 1116 118
rect 1142 114 1146 118
rect 1039 14 1043 18
rect 1069 14 1073 18
rect 1081 14 1085 18
rect 1095 14 1099 18
rect 1356 201 1360 205
rect 1651 197 1655 201
rect 1259 162 1263 166
rect 1289 162 1293 166
rect 1394 166 1398 170
rect 1424 166 1428 170
rect 1326 118 1330 122
rect 1356 118 1360 122
rect 1261 14 1265 18
rect 1291 14 1295 18
rect 1303 14 1307 18
rect 1317 14 1321 18
rect 1373 14 1377 18
rect 1387 14 1391 18
rect 1403 14 1407 18
rect 1415 14 1419 18
rect 1429 14 1433 18
rect 1681 197 1685 201
rect 1865 201 1869 205
rect 1584 158 1588 162
rect 1614 158 1618 162
rect 1719 162 1723 166
rect 1749 162 1753 166
rect 1651 114 1655 118
rect 1681 114 1685 118
rect 1578 14 1582 18
rect 1608 14 1612 18
rect 1620 14 1624 18
rect 1634 14 1638 18
rect 1895 201 1899 205
rect 1798 162 1802 166
rect 1828 162 1832 166
rect 1933 166 1937 170
rect 1963 166 1967 170
rect 1865 118 1869 122
rect 1895 118 1899 122
rect 1800 14 1804 18
rect 1830 14 1834 18
rect 1842 14 1846 18
rect 1856 14 1860 18
rect 1912 14 1916 18
rect 1926 14 1930 18
rect 1942 14 1946 18
rect 1954 14 1958 18
rect 1968 14 1972 18
<< pdcontact >>
rect 95 238 99 242
rect 110 238 114 242
rect 125 238 129 242
rect 309 242 313 246
rect 324 242 328 246
rect 339 242 343 246
rect 602 237 606 241
rect 617 237 621 241
rect 632 237 636 241
rect 816 241 820 245
rect 831 241 835 245
rect 846 241 850 245
rect 28 199 32 203
rect 43 199 47 203
rect 58 199 62 203
rect 163 203 167 207
rect 178 203 182 207
rect 193 203 197 207
rect 242 203 246 207
rect 257 203 261 207
rect 272 203 276 207
rect 95 155 99 159
rect 110 155 114 159
rect 125 155 129 159
rect 22 55 26 59
rect 37 55 41 59
rect 52 55 56 59
rect 64 55 68 59
rect 78 55 82 59
rect 377 207 381 211
rect 392 207 396 211
rect 1112 237 1116 241
rect 1127 237 1131 241
rect 1142 237 1146 241
rect 1326 241 1330 245
rect 1341 241 1345 245
rect 1356 241 1360 245
rect 407 207 411 211
rect 535 198 539 202
rect 550 198 554 202
rect 565 198 569 202
rect 309 159 313 163
rect 324 159 328 163
rect 339 159 343 163
rect 244 55 248 59
rect 259 55 263 59
rect 274 55 278 59
rect 286 55 290 59
rect 300 55 304 59
rect 356 55 360 59
rect 386 55 390 59
rect 398 55 402 59
rect 412 55 416 59
rect 670 202 674 206
rect 685 202 689 206
rect 700 202 704 206
rect 749 202 753 206
rect 764 202 768 206
rect 1651 237 1655 241
rect 1666 237 1670 241
rect 1681 237 1685 241
rect 1865 241 1869 245
rect 1880 241 1884 245
rect 1895 241 1899 245
rect 779 202 783 206
rect 602 154 606 158
rect 617 154 621 158
rect 632 154 636 158
rect 529 54 533 58
rect 544 54 548 58
rect 559 54 563 58
rect 571 54 575 58
rect 585 54 589 58
rect 884 206 888 210
rect 899 206 903 210
rect 914 206 918 210
rect 1045 198 1049 202
rect 1060 198 1064 202
rect 1075 198 1079 202
rect 816 158 820 162
rect 831 158 835 162
rect 846 158 850 162
rect 751 54 755 58
rect 766 54 770 58
rect 781 54 785 58
rect 793 54 797 58
rect 807 54 811 58
rect 863 54 867 58
rect 893 54 897 58
rect 905 54 909 58
rect 919 54 923 58
rect 1180 202 1184 206
rect 1195 202 1199 206
rect 1210 202 1214 206
rect 1259 202 1263 206
rect 1274 202 1278 206
rect 1289 202 1293 206
rect 1112 154 1116 158
rect 1127 154 1131 158
rect 1142 154 1146 158
rect 1039 54 1043 58
rect 1054 54 1058 58
rect 1069 54 1073 58
rect 1081 54 1085 58
rect 1095 54 1099 58
rect 1394 206 1398 210
rect 1409 206 1413 210
rect 1424 206 1428 210
rect 1584 198 1588 202
rect 1599 198 1603 202
rect 1614 198 1618 202
rect 1326 158 1330 162
rect 1341 158 1345 162
rect 1356 158 1360 162
rect 1261 54 1265 58
rect 1276 54 1280 58
rect 1291 54 1295 58
rect 1303 54 1307 58
rect 1317 54 1321 58
rect 1373 54 1377 58
rect 1403 54 1407 58
rect 1415 54 1419 58
rect 1429 54 1433 58
rect 1719 202 1723 206
rect 1734 202 1738 206
rect 1749 202 1753 206
rect 1798 202 1802 206
rect 1813 202 1817 206
rect 1828 202 1832 206
rect 1651 154 1655 158
rect 1666 154 1670 158
rect 1681 154 1685 158
rect 1578 54 1582 58
rect 1593 54 1597 58
rect 1608 54 1612 58
rect 1620 54 1624 58
rect 1634 54 1638 58
rect 1933 206 1937 210
rect 1948 206 1952 210
rect 1963 206 1967 210
rect 1865 158 1869 162
rect 1880 158 1884 162
rect 1895 158 1899 162
rect 1800 54 1804 58
rect 1815 54 1819 58
rect 1830 54 1834 58
rect 1842 54 1846 58
rect 1856 54 1860 58
rect 1912 54 1916 58
rect 1942 54 1946 58
rect 1954 54 1958 58
rect 1968 54 1972 58
<< nbccdiffcontact >>
rect 64 69 68 73
rect 286 69 290 73
rect 398 69 402 73
rect 571 68 575 72
rect 793 68 797 72
rect 905 68 909 72
rect 1081 68 1085 72
rect 1303 68 1307 72
rect 1415 68 1419 72
rect 1620 68 1624 72
rect 1842 68 1846 72
rect 1954 68 1958 72
<< m2contact >>
rect 303 256 307 260
rect 89 252 93 256
rect 186 252 190 256
rect 397 255 401 259
rect 61 213 65 217
rect 129 186 133 190
rect 275 217 279 221
rect 343 190 347 194
rect 810 255 814 259
rect 596 251 600 255
rect 693 251 697 255
rect 904 254 908 258
rect 63 147 67 151
rect 90 169 94 173
rect 159 151 163 155
rect 91 103 95 107
rect 129 103 133 107
rect 277 151 281 155
rect 304 173 308 177
rect 373 155 377 159
rect 305 107 309 111
rect 343 107 347 111
rect 416 76 420 80
rect 568 212 572 216
rect 636 185 640 189
rect 782 216 786 220
rect 850 189 854 193
rect 1320 255 1324 259
rect 1106 251 1110 255
rect 1203 251 1207 255
rect 1414 254 1418 258
rect 570 146 574 150
rect 597 168 601 172
rect 666 150 670 154
rect 598 102 602 106
rect 636 102 640 106
rect 784 150 788 154
rect 811 172 815 176
rect 880 154 884 158
rect 812 106 816 110
rect 850 106 854 110
rect 923 75 927 79
rect 145 5 149 9
rect 1078 212 1082 216
rect 1146 185 1150 189
rect 1292 216 1296 220
rect 1360 189 1364 193
rect 1859 255 1863 259
rect 1645 251 1649 255
rect 1742 251 1746 255
rect 1953 254 1957 258
rect 1080 146 1084 150
rect 1107 168 1111 172
rect 1176 150 1180 154
rect 1108 102 1112 106
rect 1146 102 1150 106
rect 1294 150 1298 154
rect 1321 172 1325 176
rect 1390 154 1394 158
rect 1322 106 1326 110
rect 1360 106 1364 110
rect 1433 75 1437 79
rect 1617 212 1621 216
rect 1685 185 1689 189
rect 1831 216 1835 220
rect 1899 189 1903 193
rect 1619 146 1623 150
rect 1646 168 1650 172
rect 1715 150 1719 154
rect 1647 102 1651 106
rect 1685 102 1689 106
rect 1833 150 1837 154
rect 1860 172 1864 176
rect 1929 154 1933 158
rect 1861 106 1865 110
rect 1899 106 1903 110
rect 1972 75 1976 79
rect 422 3 426 7
rect 519 2 523 7
rect 652 4 656 8
rect 925 2 929 6
rect 1035 2 1039 6
rect 1162 4 1166 8
rect 1435 2 1439 6
rect 1574 2 1578 6
rect 1701 4 1705 8
<< psubstratepcontact >>
rect 100 186 104 190
rect 121 186 125 190
rect 33 147 37 151
rect 54 147 58 151
rect 168 151 172 155
rect 189 151 193 155
rect 100 103 104 107
rect 121 103 125 107
rect 27 3 31 7
rect 48 3 52 7
rect 64 3 68 7
rect 79 3 83 7
rect 314 190 318 194
rect 335 190 339 194
rect 247 151 251 155
rect 268 151 272 155
rect 382 155 386 159
rect 403 155 407 159
rect 314 107 318 111
rect 335 107 339 111
rect 249 3 253 7
rect 270 3 274 7
rect 286 3 290 7
rect 301 3 305 7
rect 361 3 365 7
rect 382 3 386 7
rect 398 3 402 7
rect 413 3 417 7
rect 607 185 611 189
rect 628 185 632 189
rect 540 146 544 150
rect 561 146 565 150
rect 675 150 679 154
rect 696 150 700 154
rect 607 102 611 106
rect 628 102 632 106
rect 534 2 538 6
rect 555 2 559 6
rect 571 2 575 6
rect 586 2 590 6
rect 821 189 825 193
rect 842 189 846 193
rect 754 150 758 154
rect 775 150 779 154
rect 889 154 893 158
rect 910 154 914 158
rect 821 106 825 110
rect 842 106 846 110
rect 756 2 760 6
rect 777 2 781 6
rect 793 2 797 6
rect 808 2 812 6
rect 868 2 872 6
rect 889 2 893 6
rect 905 2 909 6
rect 920 2 924 6
rect 1117 185 1121 189
rect 1138 185 1142 189
rect 1050 146 1054 150
rect 1071 146 1075 150
rect 1185 150 1189 154
rect 1206 150 1210 154
rect 1117 102 1121 106
rect 1138 102 1142 106
rect 1044 2 1048 6
rect 1065 2 1069 6
rect 1081 2 1085 6
rect 1096 2 1100 6
rect 1331 189 1335 193
rect 1352 189 1356 193
rect 1264 150 1268 154
rect 1285 150 1289 154
rect 1399 154 1403 158
rect 1420 154 1424 158
rect 1331 106 1335 110
rect 1352 106 1356 110
rect 1266 2 1270 6
rect 1287 2 1291 6
rect 1303 2 1307 6
rect 1318 2 1322 6
rect 1378 2 1382 6
rect 1399 2 1403 6
rect 1415 2 1419 6
rect 1430 2 1434 6
rect 1656 185 1660 189
rect 1677 185 1681 189
rect 1589 146 1593 150
rect 1610 146 1614 150
rect 1724 150 1728 154
rect 1745 150 1749 154
rect 1656 102 1660 106
rect 1677 102 1681 106
rect 1583 2 1587 6
rect 1604 2 1608 6
rect 1620 2 1624 6
rect 1635 2 1639 6
rect 1870 189 1874 193
rect 1891 189 1895 193
rect 1803 150 1807 154
rect 1824 150 1828 154
rect 1938 154 1942 158
rect 1959 154 1963 158
rect 1870 106 1874 110
rect 1891 106 1895 110
rect 1805 2 1809 6
rect 1826 2 1830 6
rect 1842 2 1846 6
rect 1857 2 1861 6
rect 1917 2 1921 6
rect 1938 2 1942 6
rect 1954 2 1958 6
rect 1969 2 1973 6
<< nsubstratencontact >>
rect 314 256 318 260
rect 333 256 337 260
rect 100 252 104 256
rect 119 252 123 256
rect 821 255 825 259
rect 840 255 844 259
rect 1331 255 1335 259
rect 1350 255 1354 259
rect 1870 255 1874 259
rect 1889 255 1893 259
rect 607 251 611 255
rect 626 251 630 255
rect 1117 251 1121 255
rect 1136 251 1140 255
rect 1656 251 1660 255
rect 1675 251 1679 255
rect 33 213 37 217
rect 52 213 56 217
rect 168 217 172 221
rect 187 217 191 221
rect 247 217 251 221
rect 266 217 270 221
rect 382 221 386 225
rect 401 221 405 225
rect 100 169 104 173
rect 119 169 123 173
rect 27 69 31 73
rect 46 69 50 73
rect 78 69 82 73
rect 540 212 544 216
rect 559 212 563 216
rect 675 216 679 220
rect 694 216 698 220
rect 754 216 758 220
rect 773 216 777 220
rect 889 220 893 224
rect 908 220 912 224
rect 314 173 318 177
rect 333 173 337 177
rect 249 69 253 73
rect 268 69 272 73
rect 300 69 304 73
rect 361 69 365 73
rect 380 69 384 73
rect 412 69 416 73
rect 1050 212 1054 216
rect 1069 212 1073 216
rect 1185 216 1189 220
rect 1204 216 1208 220
rect 1264 216 1268 220
rect 1283 216 1287 220
rect 1399 220 1403 224
rect 1418 220 1422 224
rect 607 168 611 172
rect 626 168 630 172
rect 534 68 538 72
rect 553 68 557 72
rect 585 68 589 72
rect 821 172 825 176
rect 840 172 844 176
rect 756 68 760 72
rect 775 68 779 72
rect 807 68 811 72
rect 868 68 872 72
rect 887 68 891 72
rect 919 68 923 72
rect 1589 212 1593 216
rect 1608 212 1612 216
rect 1724 216 1728 220
rect 1743 216 1747 220
rect 1803 216 1807 220
rect 1822 216 1826 220
rect 1938 220 1942 224
rect 1957 220 1961 224
rect 1117 168 1121 172
rect 1136 168 1140 172
rect 1044 68 1048 72
rect 1063 68 1067 72
rect 1095 68 1099 72
rect 1331 172 1335 176
rect 1350 172 1354 176
rect 1266 68 1270 72
rect 1285 68 1289 72
rect 1317 68 1321 72
rect 1378 68 1382 72
rect 1397 68 1401 72
rect 1429 68 1433 72
rect 1656 168 1660 172
rect 1675 168 1679 172
rect 1583 68 1587 72
rect 1602 68 1606 72
rect 1634 68 1638 72
rect 1870 172 1874 176
rect 1889 172 1893 176
rect 1805 68 1809 72
rect 1824 68 1828 72
rect 1856 68 1860 72
rect 1917 68 1921 72
rect 1936 68 1940 72
rect 1968 68 1972 72
<< labels >>
rlabel metal1 -34 188 -34 188 3 ctrl
rlabel metal1 -15 299 -15 299 5 b3
rlabel metal1 -23 299 -23 299 5 a0
rlabel metal1 -15 299 -15 299 5 b0
rlabel metal1 484 298 484 298 5 a1
rlabel metal1 492 298 492 298 5 b1
rlabel metal1 994 298 994 298 5 a2
rlabel metal1 1002 298 1002 298 5 b2
rlabel metal1 1533 298 1533 298 5 a3
rlabel metal1 1541 298 1541 298 5 b3
rlabel polysilicon 2068 -76 2068 -76 8 s3
rlabel polysilicon 2035 -76 2035 -76 1 carry
rlabel metal1 1372 257 1372 257 1 Vdd
rlabel metal1 1356 4 1356 4 1 gnd
rlabel polysilicon 970 -76 970 -76 1 s1
rlabel polysilicon 1491 -75 1491 -75 1 s2
rlabel polysilicon 459 -75 459 -75 1 s0
<< end >>
