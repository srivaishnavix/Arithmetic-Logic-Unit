magic
tech scmos
timestamp 1701204588
<< nwell >>
rect 6 1479 133 1491
rect 896 1295 963 1307
rect 972 1295 1066 1307
rect 194 1278 292 1290
rect 301 1278 395 1290
rect 551 1280 634 1292
rect 647 1280 741 1292
rect 1302 1251 1396 1263
rect 284 1133 326 1145
rect 628 1141 670 1153
rect 986 1146 1028 1158
rect 1332 1149 1374 1161
rect 159 1094 185 1106
rect 503 1102 529 1114
rect 216 1085 258 1097
rect 351 1089 393 1101
rect 560 1093 602 1105
rect 695 1097 737 1109
rect 861 1107 887 1119
rect 918 1098 960 1110
rect 1053 1102 1095 1114
rect 1207 1110 1233 1122
rect 1264 1101 1306 1113
rect 1399 1105 1441 1117
rect 284 1050 326 1062
rect 628 1058 670 1070
rect 986 1063 1028 1075
rect 1332 1066 1374 1078
rect -99 980 -1 992
rect 1310 971 1404 983
rect 887 928 955 940
rect 964 928 1058 940
rect 180 907 278 919
rect 287 907 381 919
rect 523 915 606 927
rect 619 915 713 927
rect -47 816 80 828
rect 131 257 199 269
rect -796 196 -728 208
rect -719 196 -651 208
rect -642 196 -574 208
rect -565 196 -497 208
rect -488 196 -420 208
rect -411 196 -343 208
rect -334 196 -266 208
rect -257 196 -189 208
rect -74 181 -49 193
rect 133 181 201 193
rect 279 181 347 193
rect 449 181 517 193
rect 837 181 905 193
rect 1007 181 1075 193
rect 1342 181 1410 193
rect 1512 181 1580 193
rect 1866 181 1934 193
rect 2036 181 2104 193
rect -74 97 -49 109
rect 135 105 203 117
rect 264 67 332 79
rect 386 67 454 79
rect 556 67 624 79
rect 944 67 1012 79
rect 1114 67 1182 79
rect 1449 67 1517 79
rect 1619 67 1687 79
rect 1973 67 2041 79
rect 2143 67 2211 79
rect 137 29 205 41
rect -621 17 -553 29
rect -544 17 -476 29
rect -467 17 -399 29
rect -390 17 -322 29
rect 483 -69 525 -57
rect 996 -69 1038 -57
rect 1502 -69 1544 -57
rect 2026 -69 2068 -57
rect 416 -108 458 -96
rect 551 -104 593 -92
rect 929 -108 971 -96
rect 1064 -104 1106 -92
rect 1435 -108 1477 -96
rect 1570 -104 1612 -92
rect 1959 -108 2001 -96
rect 2094 -104 2136 -92
rect 483 -152 525 -140
rect 996 -152 1038 -140
rect 1502 -152 1544 -140
rect 2026 -152 2068 -140
rect 750 -253 792 -241
rect 985 -253 1027 -241
rect 1273 -253 1315 -241
rect 1508 -253 1550 -241
rect 1796 -253 1838 -241
rect 2031 -253 2073 -241
rect 2319 -253 2361 -241
rect 2554 -253 2596 -241
rect 683 -292 725 -280
rect 818 -288 860 -276
rect 918 -292 960 -280
rect 1053 -288 1095 -276
rect 1206 -292 1248 -280
rect 1341 -288 1383 -276
rect 1441 -292 1483 -280
rect 1576 -288 1618 -276
rect 1729 -292 1771 -280
rect 1864 -288 1906 -276
rect 1964 -292 2006 -280
rect 2099 -288 2141 -276
rect 2252 -292 2294 -280
rect 2387 -288 2429 -276
rect 2487 -292 2529 -280
rect 2622 -288 2664 -276
rect 750 -336 792 -324
rect 985 -336 1027 -324
rect 1273 -336 1315 -324
rect 1508 -336 1550 -324
rect 1796 -336 1838 -324
rect 2031 -336 2073 -324
rect 2319 -336 2361 -324
rect 2554 -336 2596 -324
rect 664 -426 732 -414
rect 916 -426 984 -414
rect 1033 -426 1101 -414
rect 1187 -426 1255 -414
rect 1439 -426 1507 -414
rect 1556 -426 1624 -414
rect 1710 -426 1778 -414
rect 1962 -426 2030 -414
rect 2079 -426 2147 -414
rect 2233 -426 2301 -414
rect 2485 -426 2553 -414
rect 2602 -426 2670 -414
<< polysilicon >>
rect 18 1530 20 1532
rect 44 1530 47 1532
rect 68 1530 71 1532
rect 94 1530 97 1532
rect 118 1530 121 1532
rect 18 1489 20 1522
rect 44 1489 47 1522
rect 68 1489 71 1522
rect 94 1489 97 1522
rect 118 1489 121 1522
rect 18 1477 20 1481
rect 44 1477 47 1481
rect 68 1477 71 1481
rect 94 1477 97 1481
rect 118 1477 121 1481
rect 136 1402 1174 1404
rect 136 1400 231 1402
rect 235 1400 588 1402
rect 592 1400 1174 1402
rect 139 1393 831 1395
rect 139 1391 246 1393
rect 250 1391 831 1393
rect 139 1381 485 1385
rect 232 1343 235 1368
rect 232 1340 240 1343
rect 237 1334 240 1340
rect 232 1331 240 1334
rect 206 1329 208 1331
rect 232 1329 235 1331
rect 247 1329 250 1368
rect 262 1329 265 1381
rect 588 1376 592 1378
rect 589 1348 592 1376
rect 589 1345 596 1348
rect 593 1335 596 1345
rect 563 1331 565 1333
rect 589 1332 596 1335
rect 589 1331 592 1332
rect 604 1331 607 1391
rect 907 1345 909 1347
rect 933 1345 936 1347
rect 948 1345 951 1347
rect 619 1331 622 1333
rect 277 1329 280 1331
rect 313 1328 315 1330
rect 339 1328 342 1330
rect 354 1328 357 1330
rect 381 1328 383 1330
rect 206 1288 208 1321
rect 232 1288 235 1321
rect 247 1288 250 1321
rect 262 1288 265 1321
rect 277 1288 280 1321
rect 659 1330 661 1332
rect 685 1330 688 1332
rect 700 1330 703 1332
rect 727 1330 729 1332
rect 313 1288 315 1320
rect 339 1307 342 1320
rect 354 1315 357 1320
rect 354 1311 358 1315
rect 339 1303 343 1307
rect 339 1288 342 1303
rect 354 1288 357 1311
rect 381 1288 383 1320
rect 397 1312 446 1316
rect 397 1295 429 1299
rect 563 1290 565 1323
rect 589 1290 592 1323
rect 604 1290 607 1323
rect 619 1290 622 1323
rect 659 1290 661 1322
rect 685 1309 688 1322
rect 700 1317 703 1322
rect 700 1313 704 1317
rect 685 1305 689 1309
rect 685 1290 688 1305
rect 700 1290 703 1313
rect 727 1290 729 1322
rect 743 1314 790 1318
rect 907 1305 909 1337
rect 933 1324 936 1337
rect 948 1332 951 1337
rect 965 1332 969 1400
rect 984 1345 986 1347
rect 1010 1345 1013 1347
rect 1025 1345 1028 1347
rect 1052 1345 1054 1347
rect 948 1328 969 1332
rect 933 1320 937 1324
rect 933 1305 936 1320
rect 948 1305 951 1328
rect 984 1305 986 1337
rect 1010 1324 1013 1337
rect 1025 1332 1028 1337
rect 1025 1328 1029 1332
rect 1010 1320 1014 1324
rect 1010 1305 1013 1320
rect 1025 1305 1028 1328
rect 1052 1305 1054 1337
rect 1068 1329 1148 1333
rect 1068 1312 1131 1316
rect 743 1297 773 1301
rect 1314 1301 1316 1303
rect 1340 1301 1343 1303
rect 1355 1301 1358 1303
rect 1382 1301 1384 1303
rect 907 1293 909 1297
rect 933 1293 936 1297
rect 948 1293 951 1297
rect 984 1293 986 1297
rect 1010 1293 1013 1297
rect 1025 1293 1028 1297
rect 1052 1293 1054 1297
rect 206 1276 208 1280
rect 232 1276 235 1280
rect 247 1276 250 1280
rect 262 1276 265 1280
rect 277 1276 280 1280
rect 313 1276 315 1280
rect 339 1276 342 1280
rect 354 1276 357 1280
rect 381 1276 383 1280
rect 563 1278 565 1282
rect 589 1278 592 1282
rect 604 1278 607 1282
rect 619 1278 622 1282
rect 659 1278 661 1282
rect 685 1278 688 1282
rect 700 1278 703 1282
rect 727 1278 729 1282
rect 1314 1261 1316 1293
rect 1340 1280 1343 1293
rect 1355 1288 1358 1293
rect 1355 1284 1359 1288
rect 1340 1276 1344 1280
rect 1340 1261 1343 1276
rect 1355 1261 1358 1284
rect 1382 1261 1384 1293
rect 1398 1285 1494 1289
rect 1398 1268 1477 1272
rect 1314 1249 1316 1253
rect 1340 1249 1343 1253
rect 1355 1249 1358 1253
rect 1382 1249 1384 1253
rect 1344 1199 1347 1201
rect 1359 1199 1362 1201
rect 998 1196 1001 1198
rect 1013 1196 1016 1198
rect 640 1191 643 1193
rect 655 1191 658 1193
rect 296 1183 299 1185
rect 311 1183 314 1185
rect 296 1162 299 1175
rect 311 1170 314 1175
rect 640 1170 643 1183
rect 655 1178 658 1183
rect 655 1174 659 1178
rect 998 1175 1001 1188
rect 1013 1183 1016 1188
rect 1013 1179 1017 1183
rect 311 1166 315 1170
rect 640 1166 644 1170
rect 296 1158 300 1162
rect 296 1143 299 1158
rect 311 1143 314 1166
rect 640 1151 643 1166
rect 655 1151 658 1174
rect 998 1171 1002 1175
rect 998 1156 1001 1171
rect 1013 1156 1016 1179
rect 1344 1178 1347 1191
rect 1359 1186 1362 1191
rect 1359 1182 1363 1186
rect 1344 1174 1348 1178
rect 1344 1159 1347 1174
rect 1359 1159 1362 1182
rect 228 1135 231 1137
rect 243 1135 246 1137
rect 363 1139 366 1141
rect 378 1139 381 1141
rect 572 1143 575 1145
rect 587 1143 590 1145
rect 707 1147 710 1149
rect 722 1147 725 1149
rect 171 1126 173 1128
rect 296 1131 299 1135
rect 311 1131 314 1135
rect 515 1134 517 1136
rect 640 1139 643 1143
rect 655 1139 658 1143
rect 930 1148 933 1150
rect 945 1148 948 1150
rect 1065 1152 1068 1154
rect 1080 1152 1083 1154
rect 873 1139 875 1141
rect 998 1144 1001 1148
rect 1013 1144 1016 1148
rect 1276 1151 1279 1153
rect 1291 1151 1294 1153
rect 1411 1155 1414 1157
rect 1426 1155 1429 1157
rect 133 1109 153 1113
rect -87 1031 -85 1033
rect -61 1031 -58 1033
rect -46 1031 -43 1033
rect -31 1031 -28 1033
rect -16 1031 -13 1033
rect 133 1028 137 1109
rect 171 1104 173 1118
rect 228 1114 231 1127
rect 243 1122 246 1127
rect 243 1118 247 1122
rect 363 1118 366 1131
rect 378 1126 381 1131
rect 378 1122 382 1126
rect 414 1122 429 1126
rect 228 1110 232 1114
rect 171 1092 173 1096
rect 228 1095 231 1110
rect 243 1095 246 1118
rect 363 1114 367 1118
rect 296 1100 299 1102
rect 311 1100 314 1102
rect 363 1099 366 1114
rect 378 1099 381 1122
rect 414 1114 446 1118
rect 515 1112 517 1126
rect 572 1122 575 1135
rect 587 1130 590 1135
rect 587 1126 591 1130
rect 707 1126 710 1139
rect 722 1134 725 1139
rect 722 1130 726 1134
rect 758 1130 773 1134
rect 572 1118 576 1122
rect 515 1100 517 1104
rect 572 1103 575 1118
rect 587 1103 590 1126
rect 707 1122 711 1126
rect 640 1108 643 1110
rect 655 1108 658 1110
rect 228 1083 231 1087
rect 243 1083 246 1087
rect 296 1079 299 1092
rect 311 1087 314 1092
rect 707 1107 710 1122
rect 722 1107 725 1130
rect 758 1122 790 1126
rect 873 1117 875 1131
rect 930 1127 933 1140
rect 945 1135 948 1140
rect 945 1131 949 1135
rect 1065 1131 1068 1144
rect 1080 1139 1083 1144
rect 1219 1142 1221 1144
rect 1344 1147 1347 1151
rect 1359 1147 1362 1151
rect 1080 1135 1084 1139
rect 1116 1135 1131 1139
rect 930 1123 934 1127
rect 572 1091 575 1095
rect 587 1091 590 1095
rect 363 1087 366 1091
rect 378 1087 381 1091
rect 640 1087 643 1100
rect 655 1095 658 1100
rect 873 1105 875 1109
rect 930 1108 933 1123
rect 945 1108 948 1131
rect 1065 1127 1069 1131
rect 998 1113 1001 1115
rect 1013 1113 1016 1115
rect 707 1095 710 1099
rect 722 1095 725 1099
rect 1065 1112 1068 1127
rect 1080 1112 1083 1135
rect 1116 1127 1148 1131
rect 1219 1120 1221 1134
rect 1276 1130 1279 1143
rect 1291 1138 1294 1143
rect 1291 1134 1295 1138
rect 1411 1134 1414 1147
rect 1426 1142 1429 1147
rect 1426 1138 1430 1142
rect 1462 1138 1477 1142
rect 1276 1126 1280 1130
rect 930 1096 933 1100
rect 945 1096 948 1100
rect 655 1091 659 1095
rect 998 1092 1001 1105
rect 1013 1100 1016 1105
rect 1219 1108 1221 1112
rect 1276 1111 1279 1126
rect 1291 1111 1294 1134
rect 1411 1130 1415 1134
rect 1344 1116 1347 1118
rect 1359 1116 1362 1118
rect 1065 1100 1068 1104
rect 1080 1100 1083 1104
rect 1411 1115 1414 1130
rect 1426 1115 1429 1138
rect 1462 1130 1494 1134
rect 1013 1096 1017 1100
rect 1276 1099 1279 1103
rect 1291 1099 1294 1103
rect 311 1083 315 1087
rect 640 1083 644 1087
rect 296 1075 300 1079
rect 296 1060 299 1075
rect 311 1060 314 1083
rect 640 1068 643 1083
rect 655 1068 658 1091
rect 998 1088 1002 1092
rect 998 1073 1001 1088
rect 1013 1073 1016 1096
rect 1344 1095 1347 1108
rect 1359 1103 1362 1108
rect 1411 1103 1414 1107
rect 1426 1103 1429 1107
rect 1359 1099 1363 1103
rect 1344 1091 1348 1095
rect 1344 1076 1347 1091
rect 1359 1076 1362 1099
rect 998 1061 1001 1065
rect 1013 1061 1016 1065
rect 1344 1064 1347 1068
rect 1359 1064 1362 1068
rect 640 1056 643 1060
rect 655 1056 658 1060
rect 296 1048 299 1052
rect 311 1048 314 1052
rect 23 1024 137 1028
rect -87 990 -85 1023
rect -61 990 -58 1023
rect -46 990 -43 1023
rect -31 990 -28 1023
rect -16 990 -13 1023
rect 23 1020 27 1024
rect 1322 1021 1324 1023
rect 1348 1021 1351 1023
rect 1363 1021 1366 1023
rect 1390 1021 1392 1023
rect 3 1016 27 1020
rect 28 1013 485 1014
rect 3 1012 485 1013
rect 3 1010 222 1012
rect 3 1009 34 1010
rect 226 1010 485 1012
rect 3 1005 34 1006
rect 3 1003 831 1005
rect 3 1002 232 1003
rect 29 1001 232 1002
rect 236 1001 564 1003
rect 568 1001 831 1003
rect 3 995 34 999
rect 30 991 1178 995
rect -87 978 -85 982
rect -61 978 -58 982
rect -46 978 -43 982
rect -31 978 -28 982
rect -16 978 -13 982
rect 223 963 226 981
rect 218 960 226 963
rect 192 958 194 960
rect 218 958 221 960
rect 233 958 236 981
rect 248 958 251 991
rect 565 970 568 979
rect 535 966 537 968
rect 561 967 568 970
rect 561 966 564 967
rect 576 966 579 991
rect 899 978 901 980
rect 925 978 928 980
rect 940 978 943 980
rect 591 966 594 968
rect 263 958 266 960
rect 299 957 301 959
rect 325 957 328 959
rect 340 957 343 959
rect 367 957 369 959
rect 631 965 633 967
rect 657 965 660 967
rect 672 965 675 967
rect 699 965 701 967
rect 192 917 194 950
rect 218 917 221 950
rect 233 917 236 950
rect 248 917 251 950
rect 263 917 266 950
rect 299 917 301 949
rect 325 936 328 949
rect 340 944 343 949
rect 340 940 344 944
rect 325 932 329 936
rect 325 917 328 932
rect 340 917 343 940
rect 367 917 369 949
rect 383 941 429 945
rect 383 924 446 928
rect 535 925 537 958
rect 561 925 564 958
rect 576 925 579 958
rect 591 925 594 958
rect 631 925 633 957
rect 657 944 660 957
rect 672 952 675 957
rect 672 948 676 952
rect 657 940 661 944
rect 657 925 660 940
rect 672 925 675 948
rect 699 925 701 957
rect 715 949 773 953
rect 899 938 901 970
rect 925 957 928 970
rect 940 965 943 970
rect 957 965 961 991
rect 1322 981 1324 1013
rect 1348 1000 1351 1013
rect 1363 1008 1366 1013
rect 1363 1004 1367 1008
rect 1348 996 1352 1000
rect 1348 981 1351 996
rect 1363 981 1366 1004
rect 1390 981 1392 1013
rect 1406 1005 1477 1009
rect 1406 988 1494 992
rect 976 978 978 980
rect 1002 978 1005 980
rect 1017 978 1020 980
rect 1044 978 1046 980
rect 940 961 961 965
rect 925 953 929 957
rect 925 938 928 953
rect 940 938 943 961
rect 976 938 978 970
rect 1002 957 1005 970
rect 1017 965 1020 970
rect 1017 961 1021 965
rect 1002 953 1006 957
rect 1002 938 1005 953
rect 1017 938 1020 961
rect 1044 938 1046 970
rect 1322 969 1324 973
rect 1348 969 1351 973
rect 1363 969 1366 973
rect 1390 969 1392 973
rect 1060 962 1131 966
rect 1060 945 1148 949
rect 715 932 790 936
rect 899 926 901 930
rect 925 926 928 930
rect 940 926 943 930
rect 976 926 978 930
rect 1002 926 1005 930
rect 1017 926 1020 930
rect 1044 926 1046 930
rect 535 913 537 917
rect 561 913 564 917
rect 576 913 579 917
rect 591 913 594 917
rect 631 913 633 917
rect 657 913 660 917
rect 672 913 675 917
rect 699 913 701 917
rect 192 905 194 909
rect 218 905 221 909
rect 233 905 236 909
rect 248 905 251 909
rect 263 905 266 909
rect 299 905 301 909
rect 325 905 328 909
rect 340 905 343 909
rect 367 905 369 909
rect -35 867 -33 869
rect -9 867 -6 869
rect 15 867 18 869
rect 41 867 44 869
rect 65 867 68 869
rect -35 826 -33 859
rect -9 826 -6 859
rect 15 826 18 859
rect 41 826 44 859
rect 65 826 68 859
rect 137 845 504 849
rect 135 838 873 842
rect 133 831 1291 835
rect -35 814 -33 818
rect -9 814 -6 818
rect 15 814 18 818
rect 41 814 44 818
rect 65 814 68 818
rect -322 576 -318 578
rect -476 476 -472 478
rect -630 371 -626 373
rect -784 311 -780 313
rect -784 206 -781 311
rect -707 296 -703 298
rect -769 206 -766 221
rect -742 206 -740 210
rect -707 206 -704 296
rect -692 206 -689 221
rect -665 206 -663 210
rect -630 206 -627 371
rect -553 352 -549 354
rect -615 206 -612 221
rect -588 206 -586 210
rect -553 206 -550 352
rect -538 206 -535 221
rect -511 206 -509 210
rect -476 206 -473 476
rect -399 462 -395 464
rect -461 206 -458 221
rect -434 206 -432 210
rect -399 206 -396 462
rect -384 206 -381 221
rect -357 206 -355 210
rect -322 206 -319 576
rect -245 537 -241 539
rect -307 206 -304 221
rect -280 206 -278 210
rect -245 206 -242 537
rect -151 331 248 335
rect -151 227 -147 331
rect 143 267 146 271
rect 158 267 161 271
rect 185 267 187 271
rect -165 223 -147 227
rect 34 240 136 244
rect -230 206 -227 221
rect -203 206 -201 210
rect -784 166 -781 198
rect -769 166 -766 198
rect -742 166 -740 198
rect -724 181 -723 185
rect -784 156 -781 158
rect -769 156 -766 158
rect -742 156 -740 158
rect -726 75 -723 181
rect -707 166 -704 198
rect -692 166 -689 198
rect -665 166 -663 198
rect -647 181 -646 185
rect -707 156 -704 158
rect -692 156 -689 158
rect -665 156 -663 158
rect -649 83 -646 181
rect -630 166 -627 198
rect -615 166 -612 198
rect -588 166 -586 198
rect -570 181 -569 185
rect -630 156 -627 158
rect -615 156 -612 158
rect -588 156 -586 158
rect -572 88 -569 181
rect -553 166 -550 198
rect -538 166 -535 198
rect -511 166 -509 198
rect -493 181 -492 185
rect -553 156 -550 158
rect -538 156 -535 158
rect -511 156 -509 158
rect -495 141 -492 181
rect -476 166 -473 198
rect -461 166 -458 198
rect -434 166 -432 198
rect -416 181 -415 185
rect -476 156 -473 158
rect -461 156 -458 158
rect -434 156 -432 158
rect -418 143 -415 181
rect -399 166 -396 198
rect -384 166 -381 198
rect -357 166 -355 198
rect -339 181 -338 185
rect -399 156 -396 158
rect -384 156 -381 158
rect -357 156 -355 158
rect -520 138 -492 141
rect -452 140 -415 143
rect -572 85 -526 88
rect -649 80 -594 83
rect -726 72 -603 75
rect -606 32 -603 72
rect -609 29 -603 32
rect -597 32 -594 80
rect -529 32 -526 85
rect -597 29 -591 32
rect -609 27 -606 29
rect -594 27 -591 29
rect -567 27 -565 31
rect -532 29 -526 32
rect -520 32 -517 138
rect -452 32 -449 140
rect -341 134 -338 181
rect -322 166 -319 198
rect -307 166 -304 198
rect -280 166 -278 198
rect -262 181 -261 185
rect -322 156 -319 158
rect -307 156 -304 158
rect -280 156 -278 158
rect -264 142 -261 181
rect -245 166 -242 198
rect -230 166 -227 198
rect -203 166 -201 198
rect -63 191 -61 195
rect -185 181 -184 185
rect -245 156 -242 158
rect -230 156 -227 158
rect -203 156 -201 158
rect -520 29 -514 32
rect -532 27 -529 29
rect -517 27 -514 29
rect -490 27 -488 31
rect -455 29 -449 32
rect -443 131 -338 134
rect -326 139 -261 142
rect -443 32 -440 131
rect -326 122 -323 139
rect -187 130 -184 181
rect -63 151 -61 183
rect -63 141 -61 143
rect -375 119 -323 122
rect -263 127 -184 130
rect 34 130 38 240
rect 143 236 146 259
rect 158 244 161 259
rect 157 240 161 244
rect -375 32 -372 119
rect -263 113 -260 127
rect 42 232 129 236
rect 142 232 146 236
rect -443 29 -437 32
rect -455 27 -452 29
rect -440 27 -437 29
rect -413 27 -411 31
rect -378 29 -372 32
rect -366 110 -260 113
rect -366 32 -363 110
rect -63 107 -61 111
rect -63 67 -61 99
rect -63 57 -61 59
rect 42 54 46 232
rect 143 227 146 232
rect 158 227 161 240
rect 185 227 187 259
rect 244 246 248 331
rect 234 242 248 246
rect 306 296 310 298
rect 143 217 146 219
rect 158 217 161 219
rect 185 217 187 219
rect 232 208 234 212
rect 145 191 148 195
rect 160 191 163 195
rect 187 191 189 195
rect 65 166 87 170
rect 83 100 87 166
rect 145 160 148 183
rect 160 168 163 183
rect 159 164 163 168
rect 144 156 148 160
rect 145 151 148 156
rect 160 151 163 164
rect 187 151 189 183
rect 232 170 236 208
rect 291 191 294 195
rect 306 191 309 296
rect 431 243 435 754
rect 413 240 435 243
rect 448 244 452 753
rect 710 336 714 338
rect 448 240 527 244
rect 413 226 416 240
rect 351 222 416 226
rect 333 191 335 195
rect 291 170 294 183
rect 234 166 294 170
rect 291 151 294 166
rect 306 151 309 183
rect 333 151 335 183
rect 351 170 355 222
rect 476 216 480 218
rect 353 166 355 170
rect 441 170 445 206
rect 461 191 464 195
rect 476 191 479 216
rect 503 191 505 195
rect 461 170 464 183
rect 441 166 464 170
rect 461 151 464 166
rect 476 151 479 183
rect 503 151 505 183
rect 523 171 527 240
rect 710 217 713 336
rect 775 225 779 754
rect 792 238 796 753
rect 1106 440 1110 442
rect 792 234 1083 238
rect 775 221 913 225
rect 710 214 867 217
rect 521 170 527 171
rect 523 166 527 170
rect 800 170 804 206
rect 849 191 852 195
rect 864 191 867 214
rect 891 191 893 195
rect 849 170 852 183
rect 800 166 852 170
rect 849 151 852 166
rect 864 151 867 183
rect 891 151 893 183
rect 909 170 913 221
rect 1034 213 1038 215
rect 911 166 913 170
rect 999 170 1003 206
rect 1019 191 1022 195
rect 1034 191 1037 213
rect 1061 191 1063 195
rect 1019 170 1022 183
rect 999 166 1022 170
rect 1019 151 1022 166
rect 1034 151 1037 183
rect 1061 151 1063 183
rect 1079 170 1083 234
rect 1106 217 1109 440
rect 1133 225 1137 753
rect 1150 238 1154 753
rect 1500 753 2112 755
rect 1496 751 2112 753
rect 1479 738 1483 751
rect 1479 734 1942 738
rect 1893 535 1897 537
rect 1150 234 1588 238
rect 1133 221 1418 225
rect 1106 214 1372 217
rect 1081 166 1083 170
rect 1305 170 1309 206
rect 1354 191 1357 195
rect 1369 191 1372 214
rect 1396 191 1398 195
rect 1354 170 1357 183
rect 1305 166 1357 170
rect 1354 151 1357 166
rect 1369 151 1372 183
rect 1396 151 1398 183
rect 1414 170 1418 221
rect 1539 213 1543 215
rect 1416 166 1418 170
rect 1504 170 1508 206
rect 1524 191 1527 195
rect 1539 191 1542 213
rect 1566 191 1568 195
rect 1524 170 1527 183
rect 1504 166 1527 170
rect 1524 151 1527 166
rect 1539 151 1542 183
rect 1566 151 1568 183
rect 1584 170 1588 234
rect 1586 166 1588 170
rect 1829 170 1833 206
rect 1878 191 1881 195
rect 1893 191 1896 535
rect 1920 191 1922 195
rect 1878 170 1881 183
rect 1829 166 1881 170
rect 1878 151 1881 166
rect 1893 151 1896 183
rect 1920 151 1922 183
rect 1938 170 1942 734
rect 2063 574 2067 576
rect 1940 166 1942 170
rect 2028 170 2032 206
rect 2048 191 2051 195
rect 2063 191 2066 574
rect 2090 191 2092 195
rect 2048 170 2051 183
rect 2028 166 2051 170
rect 2048 151 2051 166
rect 2063 151 2066 183
rect 2090 151 2092 183
rect 2108 170 2112 751
rect 2110 166 2112 170
rect 145 141 148 143
rect 160 141 163 143
rect 187 141 189 143
rect 291 141 294 143
rect 306 124 309 143
rect 333 141 335 143
rect 461 141 464 143
rect 476 141 479 143
rect 503 141 505 143
rect 849 141 852 143
rect 306 121 416 124
rect 147 115 150 119
rect 162 115 165 119
rect 189 115 191 119
rect 67 96 133 100
rect 33 50 46 54
rect -366 29 -360 32
rect -378 27 -375 29
rect -363 27 -360 29
rect -336 27 -334 31
rect -609 -13 -606 19
rect -594 -13 -591 19
rect -567 -13 -565 19
rect -551 2 -549 6
rect -609 -23 -606 -21
rect -594 -23 -591 -21
rect -567 -23 -565 -21
rect -553 -46 -549 2
rect -532 -13 -529 19
rect -517 -13 -514 19
rect -490 -13 -488 19
rect -474 2 -472 6
rect -532 -23 -529 -21
rect -517 -23 -514 -21
rect -490 -23 -488 -21
rect -476 -46 -472 2
rect -455 -13 -452 19
rect -440 -13 -437 19
rect -413 -13 -411 19
rect -397 2 -395 6
rect -455 -23 -452 -21
rect -440 -23 -437 -21
rect -413 -23 -411 -21
rect -399 -46 -395 2
rect -378 -13 -375 19
rect -363 -13 -360 19
rect -336 -13 -334 19
rect -320 2 -318 6
rect -378 -23 -375 -21
rect -363 -23 -360 -21
rect -336 -23 -334 -21
rect -322 -46 -318 2
rect 33 -213 37 50
rect 42 49 46 50
rect 58 10 62 80
rect 67 16 71 96
rect 147 84 150 107
rect 162 92 165 107
rect 161 88 165 92
rect 146 80 150 84
rect 147 75 150 80
rect 162 75 165 88
rect 189 75 191 107
rect 339 94 341 98
rect 276 77 279 81
rect 291 77 294 81
rect 318 77 320 81
rect 147 65 150 67
rect 162 65 165 67
rect 189 65 191 67
rect 276 46 279 69
rect 149 39 152 43
rect 164 39 167 43
rect 191 39 193 43
rect 275 42 279 46
rect 276 37 279 42
rect 291 37 294 69
rect 318 37 320 69
rect 339 56 343 94
rect 398 77 401 81
rect 413 77 416 121
rect 476 110 480 141
rect 864 118 867 143
rect 891 141 893 143
rect 1019 141 1022 143
rect 864 115 974 118
rect 476 106 586 110
rect 440 77 442 81
rect 398 56 401 69
rect 334 52 401 56
rect 398 37 401 52
rect 413 37 416 69
rect 440 37 442 69
rect 548 56 552 92
rect 582 89 586 106
rect 568 77 571 81
rect 583 77 586 89
rect 610 77 612 81
rect 568 56 571 69
rect 460 52 462 56
rect 548 52 571 56
rect 67 12 142 16
rect 149 8 152 31
rect 164 16 167 31
rect 163 12 167 16
rect 148 4 152 8
rect 149 -1 152 4
rect 164 -1 167 12
rect 191 -1 193 31
rect 276 27 279 29
rect 291 27 294 29
rect 318 27 320 29
rect 398 27 401 29
rect 413 27 416 29
rect 440 27 442 29
rect 458 14 462 52
rect 568 37 571 52
rect 583 37 586 69
rect 610 37 612 69
rect 907 56 911 92
rect 956 77 959 81
rect 971 77 974 115
rect 1034 116 1037 143
rect 1061 141 1063 143
rect 1354 141 1357 143
rect 1369 116 1372 143
rect 1396 141 1398 143
rect 1524 141 1527 143
rect 1539 119 1542 143
rect 1566 141 1568 143
rect 1878 141 1881 143
rect 1893 125 1896 143
rect 1920 141 1922 143
rect 2048 141 2051 143
rect 1893 122 2003 125
rect 1539 116 1649 119
rect 1034 113 1144 116
rect 1369 113 1479 116
rect 998 77 1000 81
rect 956 56 959 69
rect 630 52 632 56
rect 907 52 959 56
rect 568 27 571 29
rect 583 27 586 29
rect 610 27 612 29
rect 349 10 462 14
rect 149 -11 152 -9
rect 164 -11 167 -9
rect 191 -11 193 -9
rect 349 -121 353 10
rect 495 -59 498 -55
rect 510 -59 513 -55
rect 495 -90 498 -67
rect 510 -82 513 -67
rect 509 -86 513 -82
rect 494 -94 498 -90
rect 428 -98 431 -94
rect 443 -98 446 -94
rect 495 -99 498 -94
rect 510 -99 513 -86
rect 563 -94 566 -90
rect 578 -94 581 -90
rect 349 -125 395 -121
rect 428 -129 431 -106
rect 443 -121 446 -106
rect 495 -109 498 -107
rect 510 -109 513 -107
rect 442 -125 446 -121
rect 563 -125 566 -102
rect 578 -117 581 -102
rect 577 -121 581 -117
rect 427 -133 431 -129
rect 428 -138 431 -133
rect 443 -138 446 -125
rect 562 -129 566 -125
rect 563 -134 566 -129
rect 578 -134 581 -121
rect 495 -142 498 -138
rect 510 -142 513 -138
rect 428 -148 431 -146
rect 443 -148 446 -146
rect 563 -144 566 -142
rect 578 -144 581 -142
rect 495 -173 498 -150
rect 510 -165 513 -150
rect 509 -169 513 -165
rect 494 -177 498 -173
rect 495 -182 498 -177
rect 510 -182 513 -169
rect 495 -192 498 -190
rect 510 -192 513 -190
rect 33 -217 377 -213
rect 628 -311 632 52
rect 956 37 959 52
rect 971 37 974 69
rect 998 37 1000 69
rect 1106 56 1110 92
rect 1126 77 1129 81
rect 1141 77 1144 113
rect 1168 77 1170 81
rect 1126 56 1129 69
rect 1018 52 1020 56
rect 1106 52 1129 56
rect 956 27 959 29
rect 971 27 974 29
rect 998 27 1000 29
rect 1016 14 1020 52
rect 1126 37 1129 52
rect 1141 37 1144 69
rect 1168 37 1170 69
rect 1412 56 1416 92
rect 1461 77 1464 81
rect 1476 77 1479 113
rect 1503 77 1505 81
rect 1461 56 1464 69
rect 1188 52 1190 56
rect 1412 52 1464 56
rect 1126 27 1129 29
rect 1141 27 1144 29
rect 1168 27 1170 29
rect 907 10 1020 14
rect 907 -30 911 10
rect 1186 -25 1190 52
rect 1461 37 1464 52
rect 1476 37 1479 69
rect 1503 37 1505 69
rect 1611 56 1615 92
rect 1631 77 1634 81
rect 1646 77 1649 116
rect 1673 77 1675 81
rect 1631 56 1634 69
rect 1523 52 1525 56
rect 1611 52 1634 56
rect 1461 27 1464 29
rect 1476 27 1479 29
rect 1503 27 1505 29
rect 1521 14 1525 52
rect 1631 37 1634 52
rect 1646 37 1649 69
rect 1673 37 1675 69
rect 1936 56 1940 92
rect 1985 77 1988 81
rect 2000 77 2003 122
rect 2063 118 2066 143
rect 2090 141 2092 143
rect 2063 115 2173 118
rect 2027 77 2029 81
rect 1985 56 1988 69
rect 1693 52 1695 56
rect 1936 52 1988 56
rect 1631 27 1634 29
rect 1646 27 1649 29
rect 1673 27 1675 29
rect 1151 -29 1190 -25
rect 1412 10 1525 14
rect 636 -303 640 -123
rect 907 -121 910 -30
rect 1008 -59 1011 -55
rect 1023 -59 1026 -55
rect 1008 -90 1011 -67
rect 1023 -82 1026 -67
rect 1022 -86 1026 -82
rect 1007 -94 1011 -90
rect 941 -98 944 -94
rect 956 -98 959 -94
rect 1008 -99 1011 -94
rect 1023 -99 1026 -86
rect 1076 -94 1079 -90
rect 1091 -94 1094 -90
rect 907 -125 908 -121
rect 941 -129 944 -106
rect 956 -121 959 -106
rect 1008 -109 1011 -107
rect 1023 -109 1026 -107
rect 955 -125 959 -121
rect 1076 -125 1079 -102
rect 1091 -117 1094 -102
rect 1090 -121 1094 -117
rect 906 -133 908 -129
rect 940 -133 944 -129
rect 906 -211 910 -133
rect 941 -138 944 -133
rect 956 -138 959 -125
rect 1075 -129 1079 -125
rect 1076 -134 1079 -129
rect 1091 -134 1094 -121
rect 1008 -142 1011 -138
rect 1023 -142 1026 -138
rect 941 -148 944 -146
rect 956 -148 959 -146
rect 1076 -144 1079 -142
rect 1091 -144 1094 -142
rect 1008 -173 1011 -150
rect 1023 -165 1026 -150
rect 1022 -169 1026 -165
rect 1007 -177 1011 -173
rect 1008 -182 1011 -177
rect 1023 -182 1026 -169
rect 1008 -192 1011 -190
rect 1023 -192 1026 -190
rect 762 -243 765 -239
rect 777 -243 780 -239
rect 997 -243 1000 -239
rect 1012 -243 1015 -239
rect 762 -274 765 -251
rect 777 -266 780 -251
rect 776 -270 780 -266
rect 761 -278 765 -274
rect 695 -282 698 -278
rect 710 -282 713 -278
rect 762 -283 765 -278
rect 777 -283 780 -270
rect 997 -274 1000 -251
rect 1012 -266 1015 -251
rect 1011 -270 1015 -266
rect 830 -278 833 -274
rect 845 -278 848 -274
rect 996 -278 1000 -274
rect 654 -299 665 -296
rect 654 -410 657 -299
rect 662 -302 665 -299
rect 662 -303 666 -302
rect 695 -313 698 -290
rect 710 -305 713 -290
rect 930 -282 933 -278
rect 945 -282 948 -278
rect 762 -293 765 -291
rect 777 -293 780 -291
rect 709 -309 713 -305
rect 830 -309 833 -286
rect 845 -301 848 -286
rect 997 -283 1000 -278
rect 1012 -283 1015 -270
rect 1065 -278 1068 -274
rect 1080 -278 1083 -274
rect 844 -305 848 -301
rect 694 -317 698 -313
rect 662 -320 666 -319
rect 662 -362 665 -320
rect 695 -322 698 -317
rect 710 -322 713 -309
rect 829 -313 833 -309
rect 830 -318 833 -313
rect 845 -318 848 -305
rect 762 -326 765 -322
rect 777 -326 780 -322
rect 695 -332 698 -330
rect 710 -332 713 -330
rect 830 -328 833 -326
rect 845 -328 848 -326
rect 762 -357 765 -334
rect 777 -349 780 -334
rect 776 -353 780 -349
rect 761 -361 765 -357
rect 662 -365 687 -362
rect 684 -410 687 -365
rect 762 -366 765 -361
rect 777 -366 780 -353
rect 762 -376 765 -374
rect 777 -376 780 -374
rect 654 -413 679 -410
rect 684 -413 694 -410
rect 676 -416 679 -413
rect 691 -416 694 -413
rect 718 -416 720 -412
rect 676 -456 679 -424
rect 691 -456 694 -424
rect 718 -456 720 -424
rect 676 -466 679 -464
rect 691 -466 694 -464
rect 718 -466 720 -464
rect 734 -478 738 -437
rect 869 -447 873 -398
rect 881 -431 885 -307
rect 930 -313 933 -290
rect 945 -305 948 -290
rect 997 -293 1000 -291
rect 1012 -293 1015 -291
rect 944 -309 948 -305
rect 1065 -309 1068 -286
rect 1080 -301 1083 -286
rect 1079 -305 1083 -301
rect 929 -317 933 -313
rect 895 -390 899 -319
rect 930 -322 933 -317
rect 945 -322 948 -309
rect 1064 -313 1068 -309
rect 1065 -318 1068 -313
rect 1080 -318 1083 -305
rect 997 -326 1000 -322
rect 1012 -326 1015 -322
rect 930 -332 933 -330
rect 945 -332 948 -330
rect 1065 -328 1068 -326
rect 1080 -328 1083 -326
rect 997 -357 1000 -334
rect 1012 -349 1015 -334
rect 1011 -353 1015 -349
rect 996 -361 1000 -357
rect 997 -366 1000 -361
rect 1012 -366 1015 -353
rect 997 -376 1000 -374
rect 1012 -376 1015 -374
rect 928 -416 931 -412
rect 943 -416 946 -412
rect 970 -416 972 -412
rect 1045 -416 1048 -412
rect 1060 -416 1063 -412
rect 1087 -416 1089 -412
rect 881 -435 883 -431
rect 928 -447 931 -424
rect 943 -439 946 -424
rect 942 -443 946 -439
rect 869 -451 871 -447
rect 927 -451 931 -447
rect 928 -456 931 -451
rect 943 -456 946 -443
rect 970 -456 972 -424
rect 1045 -447 1048 -424
rect 1044 -451 1048 -447
rect 1045 -456 1048 -451
rect 1060 -456 1063 -424
rect 1087 -456 1089 -424
rect 928 -466 931 -464
rect 943 -466 946 -464
rect 970 -466 972 -464
rect 1045 -466 1048 -464
rect 1060 -466 1063 -464
rect 1087 -466 1089 -464
rect 1045 -468 1052 -466
rect 1049 -478 1052 -468
rect 734 -482 1052 -478
rect 1122 -489 1126 -307
rect 1151 -311 1155 -29
rect 1159 -303 1163 -123
rect 1412 -121 1416 10
rect 1691 -26 1695 52
rect 1985 37 1988 52
rect 2000 37 2003 69
rect 2027 37 2029 69
rect 2135 56 2139 92
rect 2155 77 2158 81
rect 2170 77 2173 115
rect 2197 77 2199 81
rect 2155 56 2158 69
rect 2047 52 2049 56
rect 2135 52 2158 56
rect 1985 27 1988 29
rect 2000 27 2003 29
rect 2027 27 2029 29
rect 2045 14 2049 52
rect 2155 37 2158 52
rect 2170 37 2173 69
rect 2197 37 2199 69
rect 2217 52 2219 56
rect 2155 27 2158 29
rect 2170 27 2173 29
rect 2197 27 2199 29
rect 1674 -30 1695 -26
rect 1936 10 2049 14
rect 1514 -59 1517 -55
rect 1529 -59 1532 -55
rect 1514 -90 1517 -67
rect 1529 -82 1532 -67
rect 1528 -86 1532 -82
rect 1513 -94 1517 -90
rect 1447 -98 1450 -94
rect 1462 -98 1465 -94
rect 1514 -99 1517 -94
rect 1529 -99 1532 -86
rect 1582 -94 1585 -90
rect 1597 -94 1600 -90
rect 1412 -125 1414 -121
rect 1447 -129 1450 -106
rect 1462 -121 1465 -106
rect 1514 -109 1517 -107
rect 1529 -109 1532 -107
rect 1461 -125 1465 -121
rect 1582 -125 1585 -102
rect 1597 -117 1600 -102
rect 1596 -121 1600 -117
rect 1412 -133 1414 -129
rect 1446 -133 1450 -129
rect 1412 -211 1416 -133
rect 1447 -138 1450 -133
rect 1462 -138 1465 -125
rect 1581 -129 1585 -125
rect 1582 -134 1585 -129
rect 1597 -134 1600 -121
rect 1514 -142 1517 -138
rect 1529 -142 1532 -138
rect 1447 -148 1450 -146
rect 1462 -148 1465 -146
rect 1582 -144 1585 -142
rect 1597 -144 1600 -142
rect 1514 -173 1517 -150
rect 1529 -165 1532 -150
rect 1528 -169 1532 -165
rect 1513 -177 1517 -173
rect 1514 -182 1517 -177
rect 1529 -182 1532 -169
rect 1514 -192 1517 -190
rect 1529 -192 1532 -190
rect 1285 -243 1288 -239
rect 1300 -243 1303 -239
rect 1520 -243 1523 -239
rect 1535 -243 1538 -239
rect 1285 -274 1288 -251
rect 1300 -266 1303 -251
rect 1299 -270 1303 -266
rect 1284 -278 1288 -274
rect 1218 -282 1221 -278
rect 1233 -282 1236 -278
rect 1285 -283 1288 -278
rect 1300 -283 1303 -270
rect 1520 -274 1523 -251
rect 1535 -266 1538 -251
rect 1534 -270 1538 -266
rect 1353 -278 1356 -274
rect 1368 -278 1371 -274
rect 1519 -278 1523 -274
rect 1177 -299 1188 -296
rect 1177 -410 1180 -299
rect 1185 -302 1188 -299
rect 1185 -303 1189 -302
rect 1218 -313 1221 -290
rect 1233 -305 1236 -290
rect 1453 -282 1456 -278
rect 1468 -282 1471 -278
rect 1285 -293 1288 -291
rect 1300 -293 1303 -291
rect 1232 -309 1236 -305
rect 1353 -309 1356 -286
rect 1368 -301 1371 -286
rect 1520 -283 1523 -278
rect 1535 -283 1538 -270
rect 1588 -278 1591 -274
rect 1603 -278 1606 -274
rect 1367 -305 1371 -301
rect 1217 -317 1221 -313
rect 1185 -320 1189 -319
rect 1185 -362 1188 -320
rect 1218 -322 1221 -317
rect 1233 -322 1236 -309
rect 1352 -313 1356 -309
rect 1353 -318 1356 -313
rect 1368 -318 1371 -305
rect 1285 -326 1288 -322
rect 1300 -326 1303 -322
rect 1218 -332 1221 -330
rect 1233 -332 1236 -330
rect 1353 -328 1356 -326
rect 1368 -328 1371 -326
rect 1285 -357 1288 -334
rect 1300 -349 1303 -334
rect 1299 -353 1303 -349
rect 1284 -361 1288 -357
rect 1185 -365 1210 -362
rect 1207 -410 1210 -365
rect 1285 -366 1288 -361
rect 1300 -366 1303 -353
rect 1285 -376 1288 -374
rect 1300 -376 1303 -374
rect 1177 -413 1202 -410
rect 1207 -413 1217 -410
rect 1199 -416 1202 -413
rect 1214 -416 1217 -413
rect 1241 -416 1243 -412
rect 1199 -456 1202 -424
rect 1214 -456 1217 -424
rect 1241 -456 1243 -424
rect 1199 -466 1202 -464
rect 1214 -466 1217 -464
rect 1241 -466 1243 -464
rect 1257 -478 1261 -437
rect 1392 -447 1396 -398
rect 1404 -431 1408 -307
rect 1453 -313 1456 -290
rect 1468 -305 1471 -290
rect 1520 -293 1523 -291
rect 1535 -293 1538 -291
rect 1467 -309 1471 -305
rect 1588 -309 1591 -286
rect 1603 -301 1606 -286
rect 1602 -305 1606 -301
rect 1452 -317 1456 -313
rect 1418 -390 1422 -319
rect 1453 -322 1456 -317
rect 1468 -322 1471 -309
rect 1587 -313 1591 -309
rect 1588 -318 1591 -313
rect 1603 -318 1606 -305
rect 1520 -326 1523 -322
rect 1535 -326 1538 -322
rect 1453 -332 1456 -330
rect 1468 -332 1471 -330
rect 1588 -328 1591 -326
rect 1603 -328 1606 -326
rect 1520 -357 1523 -334
rect 1535 -349 1538 -334
rect 1534 -353 1538 -349
rect 1519 -361 1523 -357
rect 1520 -366 1523 -361
rect 1535 -366 1538 -353
rect 1520 -376 1523 -374
rect 1535 -376 1538 -374
rect 1451 -416 1454 -412
rect 1466 -416 1469 -412
rect 1493 -416 1495 -412
rect 1568 -416 1571 -412
rect 1583 -416 1586 -412
rect 1610 -416 1612 -412
rect 1404 -435 1406 -431
rect 1451 -447 1454 -424
rect 1466 -439 1469 -424
rect 1465 -443 1469 -439
rect 1392 -451 1394 -447
rect 1450 -451 1454 -447
rect 1451 -456 1454 -451
rect 1466 -456 1469 -443
rect 1493 -456 1495 -424
rect 1568 -447 1571 -424
rect 1567 -451 1571 -447
rect 1568 -456 1571 -451
rect 1583 -456 1586 -424
rect 1610 -456 1612 -424
rect 1451 -466 1454 -464
rect 1466 -466 1469 -464
rect 1493 -466 1495 -464
rect 1568 -466 1571 -464
rect 1583 -466 1586 -464
rect 1610 -466 1612 -464
rect 1568 -468 1575 -466
rect 1572 -478 1575 -468
rect 1257 -482 1575 -478
rect 1645 -489 1649 -307
rect 1674 -311 1678 -30
rect 1682 -303 1686 -123
rect 1936 -121 1940 10
rect 2215 -26 2219 52
rect 2197 -30 2219 -26
rect 2038 -59 2041 -55
rect 2053 -59 2056 -55
rect 2038 -90 2041 -67
rect 2053 -82 2056 -67
rect 2052 -86 2056 -82
rect 2037 -94 2041 -90
rect 1971 -98 1974 -94
rect 1986 -98 1989 -94
rect 2038 -99 2041 -94
rect 2053 -99 2056 -86
rect 2106 -94 2109 -90
rect 2121 -94 2124 -90
rect 1936 -125 1938 -121
rect 1971 -129 1974 -106
rect 1986 -121 1989 -106
rect 2038 -109 2041 -107
rect 2053 -109 2056 -107
rect 1985 -125 1989 -121
rect 2106 -125 2109 -102
rect 2121 -117 2124 -102
rect 2120 -121 2124 -117
rect 1936 -133 1938 -129
rect 1970 -133 1974 -129
rect 1936 -211 1940 -133
rect 1971 -138 1974 -133
rect 1986 -138 1989 -125
rect 2105 -129 2109 -125
rect 2106 -134 2109 -129
rect 2121 -134 2124 -121
rect 2038 -142 2041 -138
rect 2053 -142 2056 -138
rect 1971 -148 1974 -146
rect 1986 -148 1989 -146
rect 2106 -144 2109 -142
rect 2121 -144 2124 -142
rect 2038 -173 2041 -150
rect 2053 -165 2056 -150
rect 2052 -169 2056 -165
rect 2037 -177 2041 -173
rect 2038 -182 2041 -177
rect 2053 -182 2056 -169
rect 2038 -192 2041 -190
rect 2053 -192 2056 -190
rect 1808 -243 1811 -239
rect 1823 -243 1826 -239
rect 2043 -243 2046 -239
rect 2058 -243 2061 -239
rect 1808 -274 1811 -251
rect 1823 -266 1826 -251
rect 1822 -270 1826 -266
rect 1807 -278 1811 -274
rect 1741 -282 1744 -278
rect 1756 -282 1759 -278
rect 1808 -283 1811 -278
rect 1823 -283 1826 -270
rect 2043 -274 2046 -251
rect 2058 -266 2061 -251
rect 2057 -270 2061 -266
rect 1876 -278 1879 -274
rect 1891 -278 1894 -274
rect 2042 -278 2046 -274
rect 1700 -299 1711 -296
rect 1700 -410 1703 -299
rect 1708 -302 1711 -299
rect 1708 -303 1712 -302
rect 1741 -313 1744 -290
rect 1756 -305 1759 -290
rect 1976 -282 1979 -278
rect 1991 -282 1994 -278
rect 1808 -293 1811 -291
rect 1823 -293 1826 -291
rect 1755 -309 1759 -305
rect 1876 -309 1879 -286
rect 1891 -301 1894 -286
rect 2043 -283 2046 -278
rect 2058 -283 2061 -270
rect 2111 -278 2114 -274
rect 2126 -278 2129 -274
rect 1890 -305 1894 -301
rect 1740 -317 1744 -313
rect 1708 -320 1712 -319
rect 1708 -362 1711 -320
rect 1741 -322 1744 -317
rect 1756 -322 1759 -309
rect 1875 -313 1879 -309
rect 1876 -318 1879 -313
rect 1891 -318 1894 -305
rect 1808 -326 1811 -322
rect 1823 -326 1826 -322
rect 1741 -332 1744 -330
rect 1756 -332 1759 -330
rect 1876 -328 1879 -326
rect 1891 -328 1894 -326
rect 1808 -357 1811 -334
rect 1823 -349 1826 -334
rect 1822 -353 1826 -349
rect 1807 -361 1811 -357
rect 1708 -365 1733 -362
rect 1730 -410 1733 -365
rect 1808 -366 1811 -361
rect 1823 -366 1826 -353
rect 1808 -376 1811 -374
rect 1823 -376 1826 -374
rect 1700 -413 1725 -410
rect 1730 -413 1740 -410
rect 1722 -416 1725 -413
rect 1737 -416 1740 -413
rect 1764 -416 1766 -412
rect 1722 -456 1725 -424
rect 1737 -456 1740 -424
rect 1764 -456 1766 -424
rect 1722 -466 1725 -464
rect 1737 -466 1740 -464
rect 1764 -466 1766 -464
rect 1780 -478 1784 -437
rect 1915 -447 1919 -398
rect 1927 -431 1931 -307
rect 1976 -313 1979 -290
rect 1991 -305 1994 -290
rect 2043 -293 2046 -291
rect 2058 -293 2061 -291
rect 1990 -309 1994 -305
rect 2111 -309 2114 -286
rect 2126 -301 2129 -286
rect 2125 -305 2129 -301
rect 1975 -317 1979 -313
rect 1941 -390 1945 -319
rect 1976 -322 1979 -317
rect 1991 -322 1994 -309
rect 2110 -313 2114 -309
rect 2111 -318 2114 -313
rect 2126 -318 2129 -305
rect 2043 -326 2046 -322
rect 2058 -326 2061 -322
rect 1976 -332 1979 -330
rect 1991 -332 1994 -330
rect 2111 -328 2114 -326
rect 2126 -328 2129 -326
rect 2043 -357 2046 -334
rect 2058 -349 2061 -334
rect 2057 -353 2061 -349
rect 2042 -361 2046 -357
rect 2043 -366 2046 -361
rect 2058 -366 2061 -353
rect 2043 -376 2046 -374
rect 2058 -376 2061 -374
rect 1974 -416 1977 -412
rect 1989 -416 1992 -412
rect 2016 -416 2018 -412
rect 2091 -416 2094 -412
rect 2106 -416 2109 -412
rect 2133 -416 2135 -412
rect 1927 -435 1929 -431
rect 1974 -447 1977 -424
rect 1989 -439 1992 -424
rect 1988 -443 1992 -439
rect 1915 -451 1917 -447
rect 1973 -451 1977 -447
rect 1974 -456 1977 -451
rect 1989 -456 1992 -443
rect 2016 -456 2018 -424
rect 2091 -447 2094 -424
rect 2090 -451 2094 -447
rect 2091 -456 2094 -451
rect 2106 -456 2109 -424
rect 2133 -456 2135 -424
rect 1974 -466 1977 -464
rect 1989 -466 1992 -464
rect 2016 -466 2018 -464
rect 2091 -466 2094 -464
rect 2106 -466 2109 -464
rect 2133 -466 2135 -464
rect 2091 -468 2098 -466
rect 2095 -478 2098 -468
rect 1780 -482 2098 -478
rect 2168 -489 2172 -307
rect 2197 -311 2201 -30
rect 2205 -303 2209 -123
rect 2331 -243 2334 -239
rect 2346 -243 2349 -239
rect 2566 -243 2569 -239
rect 2581 -243 2584 -239
rect 2331 -274 2334 -251
rect 2346 -266 2349 -251
rect 2345 -270 2349 -266
rect 2330 -278 2334 -274
rect 2264 -282 2267 -278
rect 2279 -282 2282 -278
rect 2331 -283 2334 -278
rect 2346 -283 2349 -270
rect 2566 -274 2569 -251
rect 2581 -266 2584 -251
rect 2580 -270 2584 -266
rect 2399 -278 2402 -274
rect 2414 -278 2417 -274
rect 2565 -278 2569 -274
rect 2223 -299 2234 -296
rect 2223 -410 2226 -299
rect 2231 -302 2234 -299
rect 2231 -303 2235 -302
rect 2264 -313 2267 -290
rect 2279 -305 2282 -290
rect 2499 -282 2502 -278
rect 2514 -282 2517 -278
rect 2331 -293 2334 -291
rect 2346 -293 2349 -291
rect 2278 -309 2282 -305
rect 2399 -309 2402 -286
rect 2414 -301 2417 -286
rect 2566 -283 2569 -278
rect 2581 -283 2584 -270
rect 2634 -278 2637 -274
rect 2649 -278 2652 -274
rect 2413 -305 2417 -301
rect 2263 -317 2267 -313
rect 2231 -320 2235 -319
rect 2231 -362 2234 -320
rect 2264 -322 2267 -317
rect 2279 -322 2282 -309
rect 2398 -313 2402 -309
rect 2399 -318 2402 -313
rect 2414 -318 2417 -305
rect 2331 -326 2334 -322
rect 2346 -326 2349 -322
rect 2264 -332 2267 -330
rect 2279 -332 2282 -330
rect 2399 -328 2402 -326
rect 2414 -328 2417 -326
rect 2331 -357 2334 -334
rect 2346 -349 2349 -334
rect 2345 -353 2349 -349
rect 2330 -361 2334 -357
rect 2231 -365 2256 -362
rect 2253 -410 2256 -365
rect 2331 -366 2334 -361
rect 2346 -366 2349 -353
rect 2331 -376 2334 -374
rect 2346 -376 2349 -374
rect 2223 -413 2248 -410
rect 2253 -413 2263 -410
rect 2245 -416 2248 -413
rect 2260 -416 2263 -413
rect 2287 -416 2289 -412
rect 2245 -456 2248 -424
rect 2260 -456 2263 -424
rect 2287 -456 2289 -424
rect 2245 -466 2248 -464
rect 2260 -466 2263 -464
rect 2287 -466 2289 -464
rect 2303 -478 2307 -437
rect 2438 -447 2442 -398
rect 2450 -431 2454 -307
rect 2499 -313 2502 -290
rect 2514 -305 2517 -290
rect 2566 -293 2569 -291
rect 2581 -293 2584 -291
rect 2513 -309 2517 -305
rect 2634 -309 2637 -286
rect 2649 -301 2652 -286
rect 2648 -305 2652 -301
rect 2498 -317 2502 -313
rect 2464 -390 2468 -319
rect 2499 -322 2502 -317
rect 2514 -322 2517 -309
rect 2633 -313 2637 -309
rect 2634 -318 2637 -313
rect 2649 -318 2652 -305
rect 2566 -326 2569 -322
rect 2581 -326 2584 -322
rect 2499 -332 2502 -330
rect 2514 -332 2517 -330
rect 2634 -328 2637 -326
rect 2649 -328 2652 -326
rect 2566 -357 2569 -334
rect 2581 -349 2584 -334
rect 2580 -353 2584 -349
rect 2565 -361 2569 -357
rect 2566 -366 2569 -361
rect 2581 -366 2584 -353
rect 2566 -376 2569 -374
rect 2581 -376 2584 -374
rect 2497 -416 2500 -412
rect 2512 -416 2515 -412
rect 2539 -416 2541 -412
rect 2614 -416 2617 -412
rect 2629 -416 2632 -412
rect 2656 -416 2658 -412
rect 2450 -435 2452 -431
rect 2497 -447 2500 -424
rect 2512 -439 2515 -424
rect 2511 -443 2515 -439
rect 2438 -451 2440 -447
rect 2496 -451 2500 -447
rect 2497 -456 2500 -451
rect 2512 -456 2515 -443
rect 2539 -456 2541 -424
rect 2614 -447 2617 -424
rect 2613 -451 2617 -447
rect 2614 -456 2617 -451
rect 2629 -456 2632 -424
rect 2656 -456 2658 -424
rect 2497 -466 2500 -464
rect 2512 -466 2515 -464
rect 2539 -466 2541 -464
rect 2614 -466 2617 -464
rect 2629 -466 2632 -464
rect 2656 -466 2658 -464
rect 2614 -468 2621 -466
rect 2618 -478 2621 -468
rect 2303 -482 2621 -478
rect 2691 -489 2695 -307
<< ndiffusion >>
rect 8 1528 18 1530
rect 8 1524 10 1528
rect 14 1524 18 1528
rect 8 1522 18 1524
rect 20 1528 30 1530
rect 20 1524 24 1528
rect 28 1524 30 1528
rect 20 1522 30 1524
rect 34 1528 44 1530
rect 34 1524 36 1528
rect 40 1524 44 1528
rect 34 1522 44 1524
rect 47 1528 56 1530
rect 47 1524 51 1528
rect 55 1524 56 1528
rect 47 1522 56 1524
rect 60 1528 68 1530
rect 60 1524 61 1528
rect 65 1524 68 1528
rect 60 1522 68 1524
rect 71 1528 81 1530
rect 71 1524 75 1528
rect 79 1524 81 1528
rect 71 1522 81 1524
rect 85 1528 94 1530
rect 85 1524 87 1528
rect 91 1524 94 1528
rect 85 1522 94 1524
rect 97 1528 107 1530
rect 97 1524 101 1528
rect 105 1524 107 1528
rect 97 1522 107 1524
rect 111 1528 118 1530
rect 115 1524 118 1528
rect 111 1522 118 1524
rect 121 1528 131 1530
rect 121 1524 125 1528
rect 129 1524 131 1528
rect 121 1522 131 1524
rect 897 1343 907 1345
rect 897 1339 899 1343
rect 903 1339 907 1343
rect 897 1337 907 1339
rect 909 1343 919 1345
rect 909 1339 913 1343
rect 917 1339 919 1343
rect 909 1337 919 1339
rect 923 1343 933 1345
rect 923 1339 925 1343
rect 929 1339 933 1343
rect 923 1337 933 1339
rect 936 1337 948 1345
rect 951 1343 961 1345
rect 951 1339 955 1343
rect 959 1339 961 1343
rect 951 1337 961 1339
rect 196 1327 206 1329
rect 196 1323 198 1327
rect 202 1323 206 1327
rect 196 1321 206 1323
rect 208 1327 218 1329
rect 208 1323 212 1327
rect 216 1323 218 1327
rect 208 1321 218 1323
rect 222 1327 232 1329
rect 222 1323 224 1327
rect 228 1323 232 1327
rect 222 1321 232 1323
rect 235 1321 247 1329
rect 250 1321 262 1329
rect 265 1321 277 1329
rect 280 1327 290 1329
rect 553 1329 563 1331
rect 280 1323 284 1327
rect 288 1323 290 1327
rect 280 1321 290 1323
rect 303 1326 313 1328
rect 303 1322 305 1326
rect 309 1322 313 1326
rect 303 1320 313 1322
rect 315 1326 325 1328
rect 315 1322 319 1326
rect 323 1322 325 1326
rect 315 1320 325 1322
rect 329 1326 339 1328
rect 329 1322 331 1326
rect 335 1322 339 1326
rect 329 1320 339 1322
rect 342 1320 354 1328
rect 357 1326 367 1328
rect 357 1322 361 1326
rect 365 1322 367 1326
rect 357 1320 367 1322
rect 371 1326 381 1328
rect 371 1322 373 1326
rect 377 1322 381 1326
rect 371 1320 381 1322
rect 383 1326 393 1328
rect 383 1322 387 1326
rect 391 1322 393 1326
rect 553 1325 555 1329
rect 559 1325 563 1329
rect 553 1323 563 1325
rect 565 1329 575 1331
rect 565 1325 569 1329
rect 573 1325 575 1329
rect 565 1323 575 1325
rect 579 1329 589 1331
rect 579 1325 581 1329
rect 585 1325 589 1329
rect 579 1323 589 1325
rect 592 1323 604 1331
rect 607 1323 619 1331
rect 622 1329 632 1331
rect 622 1325 626 1329
rect 630 1325 632 1329
rect 622 1323 632 1325
rect 649 1328 659 1330
rect 649 1324 651 1328
rect 655 1324 659 1328
rect 383 1320 393 1322
rect 649 1322 659 1324
rect 661 1328 671 1330
rect 661 1324 665 1328
rect 669 1324 671 1328
rect 661 1322 671 1324
rect 675 1328 685 1330
rect 675 1324 677 1328
rect 681 1324 685 1328
rect 675 1322 685 1324
rect 688 1322 700 1330
rect 703 1328 713 1330
rect 703 1324 707 1328
rect 711 1324 713 1328
rect 703 1322 713 1324
rect 717 1328 727 1330
rect 717 1324 719 1328
rect 723 1324 727 1328
rect 717 1322 727 1324
rect 729 1328 739 1330
rect 729 1324 733 1328
rect 737 1324 739 1328
rect 729 1322 739 1324
rect 974 1343 984 1345
rect 974 1339 976 1343
rect 980 1339 984 1343
rect 974 1337 984 1339
rect 986 1343 996 1345
rect 986 1339 990 1343
rect 994 1339 996 1343
rect 986 1337 996 1339
rect 1000 1343 1010 1345
rect 1000 1339 1002 1343
rect 1006 1339 1010 1343
rect 1000 1337 1010 1339
rect 1013 1337 1025 1345
rect 1028 1343 1038 1345
rect 1028 1339 1032 1343
rect 1036 1339 1038 1343
rect 1028 1337 1038 1339
rect 1042 1343 1052 1345
rect 1042 1339 1044 1343
rect 1048 1339 1052 1343
rect 1042 1337 1052 1339
rect 1054 1343 1064 1345
rect 1054 1339 1058 1343
rect 1062 1339 1064 1343
rect 1054 1337 1064 1339
rect 1304 1299 1314 1301
rect 1304 1295 1306 1299
rect 1310 1295 1314 1299
rect 1304 1293 1314 1295
rect 1316 1299 1326 1301
rect 1316 1295 1320 1299
rect 1324 1295 1326 1299
rect 1316 1293 1326 1295
rect 1330 1299 1340 1301
rect 1330 1295 1332 1299
rect 1336 1295 1340 1299
rect 1330 1293 1340 1295
rect 1343 1293 1355 1301
rect 1358 1299 1368 1301
rect 1358 1295 1362 1299
rect 1366 1295 1368 1299
rect 1358 1293 1368 1295
rect 1372 1299 1382 1301
rect 1372 1295 1374 1299
rect 1378 1295 1382 1299
rect 1372 1293 1382 1295
rect 1384 1299 1394 1301
rect 1384 1295 1388 1299
rect 1392 1295 1394 1299
rect 1384 1293 1394 1295
rect 1334 1197 1344 1199
rect 988 1194 998 1196
rect 630 1189 640 1191
rect 630 1185 632 1189
rect 636 1185 640 1189
rect 630 1183 640 1185
rect 643 1183 655 1191
rect 658 1189 668 1191
rect 658 1185 662 1189
rect 666 1185 668 1189
rect 988 1190 990 1194
rect 994 1190 998 1194
rect 988 1188 998 1190
rect 1001 1188 1013 1196
rect 1016 1194 1026 1196
rect 1016 1190 1020 1194
rect 1024 1190 1026 1194
rect 1334 1193 1336 1197
rect 1340 1193 1344 1197
rect 1334 1191 1344 1193
rect 1347 1191 1359 1199
rect 1362 1197 1372 1199
rect 1362 1193 1366 1197
rect 1370 1193 1372 1197
rect 1362 1191 1372 1193
rect 1016 1188 1026 1190
rect 658 1183 668 1185
rect 286 1181 296 1183
rect 286 1177 288 1181
rect 292 1177 296 1181
rect 286 1175 296 1177
rect 299 1175 311 1183
rect 314 1181 324 1183
rect 314 1177 318 1181
rect 322 1177 324 1181
rect 314 1175 324 1177
rect 697 1145 707 1147
rect 562 1141 572 1143
rect 353 1137 363 1139
rect 218 1133 228 1135
rect 218 1129 220 1133
rect 224 1129 228 1133
rect 218 1127 228 1129
rect 231 1127 243 1135
rect 246 1133 256 1135
rect 246 1129 250 1133
rect 254 1129 256 1133
rect 353 1133 355 1137
rect 359 1133 363 1137
rect 353 1131 363 1133
rect 366 1131 378 1139
rect 381 1137 391 1139
rect 381 1133 385 1137
rect 389 1133 391 1137
rect 562 1137 564 1141
rect 568 1137 572 1141
rect 562 1135 572 1137
rect 575 1135 587 1143
rect 590 1141 600 1143
rect 590 1137 594 1141
rect 598 1137 600 1141
rect 697 1141 699 1145
rect 703 1141 707 1145
rect 697 1139 707 1141
rect 710 1139 722 1147
rect 725 1145 735 1147
rect 1055 1150 1065 1152
rect 920 1146 930 1148
rect 725 1141 729 1145
rect 733 1141 735 1145
rect 920 1142 922 1146
rect 926 1142 930 1146
rect 725 1139 735 1141
rect 920 1140 930 1142
rect 933 1140 945 1148
rect 948 1146 958 1148
rect 948 1142 952 1146
rect 956 1142 958 1146
rect 1055 1146 1057 1150
rect 1061 1146 1065 1150
rect 1055 1144 1065 1146
rect 1068 1144 1080 1152
rect 1083 1150 1093 1152
rect 1083 1146 1087 1150
rect 1091 1146 1093 1150
rect 1401 1153 1411 1155
rect 1266 1149 1276 1151
rect 1083 1144 1093 1146
rect 1266 1145 1268 1149
rect 1272 1145 1276 1149
rect 948 1140 958 1142
rect 590 1135 600 1137
rect 381 1131 391 1133
rect 505 1132 515 1134
rect 246 1127 256 1129
rect 161 1124 171 1126
rect 161 1120 163 1124
rect 167 1120 171 1124
rect 161 1118 171 1120
rect 173 1124 183 1126
rect 173 1120 177 1124
rect 181 1120 183 1124
rect 173 1118 183 1120
rect -97 1029 -87 1031
rect -97 1025 -95 1029
rect -91 1025 -87 1029
rect -97 1023 -87 1025
rect -85 1029 -75 1031
rect -85 1025 -81 1029
rect -77 1025 -75 1029
rect -85 1023 -75 1025
rect -71 1029 -61 1031
rect -71 1025 -69 1029
rect -65 1025 -61 1029
rect -71 1023 -61 1025
rect -58 1023 -46 1031
rect -43 1023 -31 1031
rect -28 1023 -16 1031
rect -13 1029 -3 1031
rect -13 1025 -9 1029
rect -5 1025 -3 1029
rect 505 1128 507 1132
rect 511 1128 515 1132
rect 505 1126 515 1128
rect 517 1132 527 1134
rect 517 1128 521 1132
rect 525 1128 527 1132
rect 517 1126 527 1128
rect 286 1098 296 1100
rect 286 1094 288 1098
rect 292 1094 296 1098
rect 286 1092 296 1094
rect 299 1092 311 1100
rect 314 1098 324 1100
rect 863 1137 873 1139
rect 863 1133 865 1137
rect 869 1133 873 1137
rect 863 1131 873 1133
rect 875 1137 885 1139
rect 875 1133 879 1137
rect 883 1133 885 1137
rect 875 1131 885 1133
rect 630 1106 640 1108
rect 314 1094 318 1098
rect 322 1094 324 1098
rect 314 1092 324 1094
rect 630 1102 632 1106
rect 636 1102 640 1106
rect 630 1100 640 1102
rect 643 1100 655 1108
rect 658 1106 668 1108
rect 1266 1143 1276 1145
rect 1279 1143 1291 1151
rect 1294 1149 1304 1151
rect 1294 1145 1298 1149
rect 1302 1145 1304 1149
rect 1401 1149 1403 1153
rect 1407 1149 1411 1153
rect 1401 1147 1411 1149
rect 1414 1147 1426 1155
rect 1429 1153 1439 1155
rect 1429 1149 1433 1153
rect 1437 1149 1439 1153
rect 1429 1147 1439 1149
rect 1294 1143 1304 1145
rect 1209 1140 1219 1142
rect 1209 1136 1211 1140
rect 1215 1136 1219 1140
rect 658 1102 662 1106
rect 666 1102 668 1106
rect 658 1100 668 1102
rect 988 1111 998 1113
rect 988 1107 990 1111
rect 994 1107 998 1111
rect 988 1105 998 1107
rect 1001 1105 1013 1113
rect 1016 1111 1026 1113
rect 1209 1134 1219 1136
rect 1221 1140 1231 1142
rect 1221 1136 1225 1140
rect 1229 1136 1231 1140
rect 1221 1134 1231 1136
rect 1016 1107 1020 1111
rect 1024 1107 1026 1111
rect 1016 1105 1026 1107
rect 1334 1114 1344 1116
rect 1334 1110 1336 1114
rect 1340 1110 1344 1114
rect 1334 1108 1344 1110
rect 1347 1108 1359 1116
rect 1362 1114 1372 1116
rect 1362 1110 1366 1114
rect 1370 1110 1372 1114
rect 1362 1108 1372 1110
rect -13 1023 -3 1025
rect 1312 1019 1322 1021
rect 1312 1015 1314 1019
rect 1318 1015 1322 1019
rect 1312 1013 1322 1015
rect 1324 1019 1334 1021
rect 1324 1015 1328 1019
rect 1332 1015 1334 1019
rect 1324 1013 1334 1015
rect 1338 1019 1348 1021
rect 1338 1015 1340 1019
rect 1344 1015 1348 1019
rect 1338 1013 1348 1015
rect 1351 1013 1363 1021
rect 1366 1019 1376 1021
rect 1366 1015 1370 1019
rect 1374 1015 1376 1019
rect 1366 1013 1376 1015
rect 1380 1019 1390 1021
rect 1380 1015 1382 1019
rect 1386 1015 1390 1019
rect 1380 1013 1390 1015
rect 1392 1019 1402 1021
rect 1392 1015 1396 1019
rect 1400 1015 1402 1019
rect 1392 1013 1402 1015
rect 889 976 899 978
rect 889 972 891 976
rect 895 972 899 976
rect 889 970 899 972
rect 901 976 911 978
rect 901 972 905 976
rect 909 972 911 976
rect 901 970 911 972
rect 915 976 925 978
rect 915 972 917 976
rect 921 972 925 976
rect 915 970 925 972
rect 928 970 940 978
rect 943 976 953 978
rect 943 972 947 976
rect 951 972 953 976
rect 943 970 953 972
rect 525 964 535 966
rect 525 960 527 964
rect 531 960 535 964
rect 182 956 192 958
rect 182 952 184 956
rect 188 952 192 956
rect 182 950 192 952
rect 194 956 204 958
rect 194 952 198 956
rect 202 952 204 956
rect 194 950 204 952
rect 208 956 218 958
rect 208 952 210 956
rect 214 952 218 956
rect 208 950 218 952
rect 221 950 233 958
rect 236 950 248 958
rect 251 950 263 958
rect 266 956 276 958
rect 525 958 535 960
rect 537 964 547 966
rect 537 960 541 964
rect 545 960 547 964
rect 537 958 547 960
rect 551 964 561 966
rect 551 960 553 964
rect 557 960 561 964
rect 551 958 561 960
rect 564 958 576 966
rect 579 958 591 966
rect 594 964 604 966
rect 594 960 598 964
rect 602 960 604 964
rect 594 958 604 960
rect 621 963 631 965
rect 621 959 623 963
rect 627 959 631 963
rect 266 952 270 956
rect 274 952 276 956
rect 266 950 276 952
rect 289 955 299 957
rect 289 951 291 955
rect 295 951 299 955
rect 289 949 299 951
rect 301 955 311 957
rect 301 951 305 955
rect 309 951 311 955
rect 301 949 311 951
rect 315 955 325 957
rect 315 951 317 955
rect 321 951 325 955
rect 315 949 325 951
rect 328 949 340 957
rect 343 955 353 957
rect 343 951 347 955
rect 351 951 353 955
rect 343 949 353 951
rect 357 955 367 957
rect 357 951 359 955
rect 363 951 367 955
rect 357 949 367 951
rect 369 955 379 957
rect 369 951 373 955
rect 377 951 379 955
rect 369 949 379 951
rect 621 957 631 959
rect 633 963 643 965
rect 633 959 637 963
rect 641 959 643 963
rect 633 957 643 959
rect 647 963 657 965
rect 647 959 649 963
rect 653 959 657 963
rect 647 957 657 959
rect 660 957 672 965
rect 675 963 685 965
rect 675 959 679 963
rect 683 959 685 963
rect 675 957 685 959
rect 689 963 699 965
rect 689 959 691 963
rect 695 959 699 963
rect 689 957 699 959
rect 701 963 711 965
rect 701 959 705 963
rect 709 959 711 963
rect 701 957 711 959
rect 966 976 976 978
rect 966 972 968 976
rect 972 972 976 976
rect 966 970 976 972
rect 978 976 988 978
rect 978 972 982 976
rect 986 972 988 976
rect 978 970 988 972
rect 992 976 1002 978
rect 992 972 994 976
rect 998 972 1002 976
rect 992 970 1002 972
rect 1005 970 1017 978
rect 1020 976 1030 978
rect 1020 972 1024 976
rect 1028 972 1030 976
rect 1020 970 1030 972
rect 1034 976 1044 978
rect 1034 972 1036 976
rect 1040 972 1044 976
rect 1034 970 1044 972
rect 1046 976 1056 978
rect 1046 972 1050 976
rect 1054 972 1056 976
rect 1046 970 1056 972
rect -45 865 -35 867
rect -45 861 -43 865
rect -39 861 -35 865
rect -45 859 -35 861
rect -33 865 -23 867
rect -33 861 -29 865
rect -25 861 -23 865
rect -33 859 -23 861
rect -19 865 -9 867
rect -19 861 -17 865
rect -13 861 -9 865
rect -19 859 -9 861
rect -6 865 3 867
rect -6 861 -2 865
rect 2 861 3 865
rect -6 859 3 861
rect 7 865 15 867
rect 7 861 8 865
rect 12 861 15 865
rect 7 859 15 861
rect 18 865 28 867
rect 18 861 22 865
rect 26 861 28 865
rect 18 859 28 861
rect 32 865 41 867
rect 32 861 34 865
rect 38 861 41 865
rect 32 859 41 861
rect 44 865 54 867
rect 44 861 48 865
rect 52 861 54 865
rect 44 859 54 861
rect 58 865 65 867
rect 62 861 65 865
rect 58 859 65 861
rect 68 865 78 867
rect 68 861 72 865
rect 76 861 78 865
rect 68 859 78 861
rect -794 164 -784 166
rect -794 160 -792 164
rect -788 160 -784 164
rect -794 158 -784 160
rect -781 158 -769 166
rect -766 164 -756 166
rect -766 160 -762 164
rect -758 160 -756 164
rect -766 158 -756 160
rect -752 164 -742 166
rect -752 160 -750 164
rect -746 160 -742 164
rect -752 158 -742 160
rect -740 164 -730 166
rect -740 160 -736 164
rect -732 160 -730 164
rect -740 158 -730 160
rect -717 164 -707 166
rect -717 160 -715 164
rect -711 160 -707 164
rect -717 158 -707 160
rect -704 158 -692 166
rect -689 164 -679 166
rect -689 160 -685 164
rect -681 160 -679 164
rect -689 158 -679 160
rect -675 164 -665 166
rect -675 160 -673 164
rect -669 160 -665 164
rect -675 158 -665 160
rect -663 164 -653 166
rect -663 160 -659 164
rect -655 160 -653 164
rect -663 158 -653 160
rect -640 164 -630 166
rect -640 160 -638 164
rect -634 160 -630 164
rect -640 158 -630 160
rect -627 158 -615 166
rect -612 164 -602 166
rect -612 160 -608 164
rect -604 160 -602 164
rect -612 158 -602 160
rect -598 164 -588 166
rect -598 160 -596 164
rect -592 160 -588 164
rect -598 158 -588 160
rect -586 164 -576 166
rect -586 160 -582 164
rect -578 160 -576 164
rect -586 158 -576 160
rect -563 164 -553 166
rect -563 160 -561 164
rect -557 160 -553 164
rect -563 158 -553 160
rect -550 158 -538 166
rect -535 164 -525 166
rect -535 160 -531 164
rect -527 160 -525 164
rect -535 158 -525 160
rect -521 164 -511 166
rect -521 160 -519 164
rect -515 160 -511 164
rect -521 158 -511 160
rect -509 164 -499 166
rect -509 160 -505 164
rect -501 160 -499 164
rect -509 158 -499 160
rect -486 164 -476 166
rect -486 160 -484 164
rect -480 160 -476 164
rect -486 158 -476 160
rect -473 158 -461 166
rect -458 164 -448 166
rect -458 160 -454 164
rect -450 160 -448 164
rect -458 158 -448 160
rect -444 164 -434 166
rect -444 160 -442 164
rect -438 160 -434 164
rect -444 158 -434 160
rect -432 164 -422 166
rect -432 160 -428 164
rect -424 160 -422 164
rect -432 158 -422 160
rect -409 164 -399 166
rect -409 160 -407 164
rect -403 160 -399 164
rect -409 158 -399 160
rect -396 158 -384 166
rect -381 164 -371 166
rect -381 160 -377 164
rect -373 160 -371 164
rect -381 158 -371 160
rect -367 164 -357 166
rect -367 160 -365 164
rect -361 160 -357 164
rect -367 158 -357 160
rect -355 164 -345 166
rect -355 160 -351 164
rect -347 160 -345 164
rect -355 158 -345 160
rect -332 164 -322 166
rect -332 160 -330 164
rect -326 160 -322 164
rect -332 158 -322 160
rect -319 158 -307 166
rect -304 164 -294 166
rect -304 160 -300 164
rect -296 160 -294 164
rect -304 158 -294 160
rect -290 164 -280 166
rect -290 160 -288 164
rect -284 160 -280 164
rect -290 158 -280 160
rect -278 164 -268 166
rect -278 160 -274 164
rect -270 160 -268 164
rect -278 158 -268 160
rect -255 164 -245 166
rect -255 160 -253 164
rect -249 160 -245 164
rect -255 158 -245 160
rect -242 158 -230 166
rect -227 164 -217 166
rect -227 160 -223 164
rect -219 160 -217 164
rect -227 158 -217 160
rect -213 164 -203 166
rect -213 160 -211 164
rect -207 160 -203 164
rect -213 158 -203 160
rect -201 164 -191 166
rect -201 160 -197 164
rect -193 160 -191 164
rect -201 158 -191 160
rect -73 149 -63 151
rect -73 145 -71 149
rect -67 145 -63 149
rect -73 143 -63 145
rect -61 149 -51 151
rect -61 145 -57 149
rect -53 145 -51 149
rect -61 143 -51 145
rect -73 65 -63 67
rect -73 61 -71 65
rect -67 61 -63 65
rect -73 59 -63 61
rect -61 65 -51 67
rect -61 61 -57 65
rect -53 61 -51 65
rect -61 59 -51 61
rect 133 225 143 227
rect 133 221 135 225
rect 139 221 143 225
rect 133 219 143 221
rect 146 219 158 227
rect 161 225 171 227
rect 161 221 165 225
rect 169 221 171 225
rect 161 219 171 221
rect 175 225 185 227
rect 175 221 177 225
rect 181 221 185 225
rect 175 219 185 221
rect 187 225 197 227
rect 187 221 191 225
rect 195 221 197 225
rect 187 219 197 221
rect 135 149 145 151
rect 135 145 137 149
rect 141 145 145 149
rect 135 143 145 145
rect 148 143 160 151
rect 163 149 173 151
rect 163 145 167 149
rect 171 145 173 149
rect 163 143 173 145
rect 177 149 187 151
rect 177 145 179 149
rect 183 145 187 149
rect 177 143 187 145
rect 189 149 199 151
rect 189 145 193 149
rect 197 145 199 149
rect 189 143 199 145
rect 281 149 291 151
rect 281 145 283 149
rect 287 145 291 149
rect 281 143 291 145
rect 294 143 306 151
rect 309 149 319 151
rect 309 145 313 149
rect 317 145 319 149
rect 309 143 319 145
rect 323 149 333 151
rect 323 145 325 149
rect 329 145 333 149
rect 323 143 333 145
rect 335 149 345 151
rect 335 145 339 149
rect 343 145 345 149
rect 335 143 345 145
rect 451 149 461 151
rect 451 145 453 149
rect 457 145 461 149
rect 451 143 461 145
rect 464 143 476 151
rect 479 149 489 151
rect 479 145 483 149
rect 487 145 489 149
rect 479 143 489 145
rect 493 149 503 151
rect 493 145 495 149
rect 499 145 503 149
rect 493 143 503 145
rect 505 149 515 151
rect 505 145 509 149
rect 513 145 515 149
rect 505 143 515 145
rect 839 149 849 151
rect 839 145 841 149
rect 845 145 849 149
rect 839 143 849 145
rect 852 143 864 151
rect 867 149 877 151
rect 867 145 871 149
rect 875 145 877 149
rect 867 143 877 145
rect 881 149 891 151
rect 881 145 883 149
rect 887 145 891 149
rect 881 143 891 145
rect 893 149 903 151
rect 893 145 897 149
rect 901 145 903 149
rect 893 143 903 145
rect 1009 149 1019 151
rect 1009 145 1011 149
rect 1015 145 1019 149
rect 1009 143 1019 145
rect 1022 143 1034 151
rect 1037 149 1047 151
rect 1037 145 1041 149
rect 1045 145 1047 149
rect 1037 143 1047 145
rect 1051 149 1061 151
rect 1051 145 1053 149
rect 1057 145 1061 149
rect 1051 143 1061 145
rect 1063 149 1073 151
rect 1063 145 1067 149
rect 1071 145 1073 149
rect 1063 143 1073 145
rect 1344 149 1354 151
rect 1344 145 1346 149
rect 1350 145 1354 149
rect 1344 143 1354 145
rect 1357 143 1369 151
rect 1372 149 1382 151
rect 1372 145 1376 149
rect 1380 145 1382 149
rect 1372 143 1382 145
rect 1386 149 1396 151
rect 1386 145 1388 149
rect 1392 145 1396 149
rect 1386 143 1396 145
rect 1398 149 1408 151
rect 1398 145 1402 149
rect 1406 145 1408 149
rect 1398 143 1408 145
rect 1514 149 1524 151
rect 1514 145 1516 149
rect 1520 145 1524 149
rect 1514 143 1524 145
rect 1527 143 1539 151
rect 1542 149 1552 151
rect 1542 145 1546 149
rect 1550 145 1552 149
rect 1542 143 1552 145
rect 1556 149 1566 151
rect 1556 145 1558 149
rect 1562 145 1566 149
rect 1556 143 1566 145
rect 1568 149 1578 151
rect 1568 145 1572 149
rect 1576 145 1578 149
rect 1568 143 1578 145
rect 1868 149 1878 151
rect 1868 145 1870 149
rect 1874 145 1878 149
rect 1868 143 1878 145
rect 1881 143 1893 151
rect 1896 149 1906 151
rect 1896 145 1900 149
rect 1904 145 1906 149
rect 1896 143 1906 145
rect 1910 149 1920 151
rect 1910 145 1912 149
rect 1916 145 1920 149
rect 1910 143 1920 145
rect 1922 149 1932 151
rect 1922 145 1926 149
rect 1930 145 1932 149
rect 1922 143 1932 145
rect 2038 149 2048 151
rect 2038 145 2040 149
rect 2044 145 2048 149
rect 2038 143 2048 145
rect 2051 143 2063 151
rect 2066 149 2076 151
rect 2066 145 2070 149
rect 2074 145 2076 149
rect 2066 143 2076 145
rect 2080 149 2090 151
rect 2080 145 2082 149
rect 2086 145 2090 149
rect 2080 143 2090 145
rect 2092 149 2102 151
rect 2092 145 2096 149
rect 2100 145 2102 149
rect 2092 143 2102 145
rect -619 -15 -609 -13
rect -619 -19 -617 -15
rect -613 -19 -609 -15
rect -619 -21 -609 -19
rect -606 -21 -594 -13
rect -591 -15 -581 -13
rect -591 -19 -587 -15
rect -583 -19 -581 -15
rect -591 -21 -581 -19
rect -577 -15 -567 -13
rect -577 -19 -575 -15
rect -571 -19 -567 -15
rect -577 -21 -567 -19
rect -565 -15 -555 -13
rect -565 -19 -561 -15
rect -557 -19 -555 -15
rect -565 -21 -555 -19
rect -542 -15 -532 -13
rect -542 -19 -540 -15
rect -536 -19 -532 -15
rect -542 -21 -532 -19
rect -529 -21 -517 -13
rect -514 -15 -504 -13
rect -514 -19 -510 -15
rect -506 -19 -504 -15
rect -514 -21 -504 -19
rect -500 -15 -490 -13
rect -500 -19 -498 -15
rect -494 -19 -490 -15
rect -500 -21 -490 -19
rect -488 -15 -478 -13
rect -488 -19 -484 -15
rect -480 -19 -478 -15
rect -488 -21 -478 -19
rect -465 -15 -455 -13
rect -465 -19 -463 -15
rect -459 -19 -455 -15
rect -465 -21 -455 -19
rect -452 -21 -440 -13
rect -437 -15 -427 -13
rect -437 -19 -433 -15
rect -429 -19 -427 -15
rect -437 -21 -427 -19
rect -423 -15 -413 -13
rect -423 -19 -421 -15
rect -417 -19 -413 -15
rect -423 -21 -413 -19
rect -411 -15 -401 -13
rect -411 -19 -407 -15
rect -403 -19 -401 -15
rect -411 -21 -401 -19
rect -388 -15 -378 -13
rect -388 -19 -386 -15
rect -382 -19 -378 -15
rect -388 -21 -378 -19
rect -375 -21 -363 -13
rect -360 -15 -350 -13
rect -360 -19 -356 -15
rect -352 -19 -350 -15
rect -360 -21 -350 -19
rect -346 -15 -336 -13
rect -346 -19 -344 -15
rect -340 -19 -336 -15
rect -346 -21 -336 -19
rect -334 -15 -324 -13
rect -334 -19 -330 -15
rect -326 -19 -324 -15
rect -334 -21 -324 -19
rect 137 73 147 75
rect 137 69 139 73
rect 143 69 147 73
rect 137 67 147 69
rect 150 67 162 75
rect 165 73 175 75
rect 165 69 169 73
rect 173 69 175 73
rect 165 67 175 69
rect 179 73 189 75
rect 179 69 181 73
rect 185 69 189 73
rect 179 67 189 69
rect 191 73 201 75
rect 191 69 195 73
rect 199 69 201 73
rect 191 67 201 69
rect 266 35 276 37
rect 266 31 268 35
rect 272 31 276 35
rect 266 29 276 31
rect 279 35 291 37
rect 279 31 282 35
rect 286 31 291 35
rect 279 29 291 31
rect 294 35 304 37
rect 294 31 298 35
rect 302 31 304 35
rect 294 29 304 31
rect 308 35 318 37
rect 308 31 310 35
rect 314 31 318 35
rect 308 29 318 31
rect 320 35 330 37
rect 320 31 324 35
rect 328 31 330 35
rect 320 29 330 31
rect 388 35 398 37
rect 388 31 390 35
rect 394 31 398 35
rect 388 29 398 31
rect 401 29 413 37
rect 416 35 426 37
rect 416 31 420 35
rect 424 31 426 35
rect 416 29 426 31
rect 430 35 440 37
rect 430 31 432 35
rect 436 31 440 35
rect 430 29 440 31
rect 442 35 452 37
rect 442 31 446 35
rect 450 31 452 35
rect 442 29 452 31
rect 558 35 568 37
rect 558 31 560 35
rect 564 31 568 35
rect 558 29 568 31
rect 571 29 583 37
rect 586 35 596 37
rect 586 31 590 35
rect 594 31 596 35
rect 586 29 596 31
rect 600 35 610 37
rect 600 31 602 35
rect 606 31 610 35
rect 600 29 610 31
rect 612 35 622 37
rect 612 31 616 35
rect 620 31 622 35
rect 612 29 622 31
rect 139 -3 149 -1
rect 139 -7 141 -3
rect 145 -7 149 -3
rect 139 -9 149 -7
rect 152 -9 164 -1
rect 167 -3 177 -1
rect 167 -7 171 -3
rect 175 -7 177 -3
rect 167 -9 177 -7
rect 181 -3 191 -1
rect 181 -7 183 -3
rect 187 -7 191 -3
rect 181 -9 191 -7
rect 193 -3 203 -1
rect 193 -7 197 -3
rect 201 -7 203 -3
rect 193 -9 203 -7
rect 485 -101 495 -99
rect 485 -105 487 -101
rect 491 -105 495 -101
rect 485 -107 495 -105
rect 498 -107 510 -99
rect 513 -101 523 -99
rect 513 -105 517 -101
rect 521 -105 523 -101
rect 513 -107 523 -105
rect 553 -136 563 -134
rect 418 -140 428 -138
rect 418 -144 420 -140
rect 424 -144 428 -140
rect 418 -146 428 -144
rect 431 -146 443 -138
rect 446 -140 456 -138
rect 446 -144 450 -140
rect 454 -144 456 -140
rect 553 -140 555 -136
rect 559 -140 563 -136
rect 553 -142 563 -140
rect 566 -142 578 -134
rect 581 -136 591 -134
rect 581 -140 585 -136
rect 589 -140 591 -136
rect 581 -142 591 -140
rect 446 -146 456 -144
rect 485 -184 495 -182
rect 485 -188 487 -184
rect 491 -188 495 -184
rect 485 -190 495 -188
rect 498 -190 510 -182
rect 513 -184 523 -182
rect 513 -188 517 -184
rect 521 -188 523 -184
rect 513 -190 523 -188
rect 946 35 956 37
rect 946 31 948 35
rect 952 31 956 35
rect 946 29 956 31
rect 959 29 971 37
rect 974 35 984 37
rect 974 31 978 35
rect 982 31 984 35
rect 974 29 984 31
rect 988 35 998 37
rect 988 31 990 35
rect 994 31 998 35
rect 988 29 998 31
rect 1000 35 1010 37
rect 1000 31 1004 35
rect 1008 31 1010 35
rect 1000 29 1010 31
rect 1116 35 1126 37
rect 1116 31 1118 35
rect 1122 31 1126 35
rect 1116 29 1126 31
rect 1129 29 1141 37
rect 1144 35 1154 37
rect 1144 31 1148 35
rect 1152 31 1154 35
rect 1144 29 1154 31
rect 1158 35 1168 37
rect 1158 31 1160 35
rect 1164 31 1168 35
rect 1158 29 1168 31
rect 1170 35 1180 37
rect 1170 31 1174 35
rect 1178 31 1180 35
rect 1170 29 1180 31
rect 1451 35 1461 37
rect 1451 31 1453 35
rect 1457 31 1461 35
rect 1451 29 1461 31
rect 1464 29 1476 37
rect 1479 35 1489 37
rect 1479 31 1483 35
rect 1487 31 1489 35
rect 1479 29 1489 31
rect 1493 35 1503 37
rect 1493 31 1495 35
rect 1499 31 1503 35
rect 1493 29 1503 31
rect 1505 35 1515 37
rect 1505 31 1509 35
rect 1513 31 1515 35
rect 1505 29 1515 31
rect 1621 35 1631 37
rect 1621 31 1623 35
rect 1627 31 1631 35
rect 1621 29 1631 31
rect 1634 29 1646 37
rect 1649 35 1659 37
rect 1649 31 1653 35
rect 1657 31 1659 35
rect 1649 29 1659 31
rect 1663 35 1673 37
rect 1663 31 1665 35
rect 1669 31 1673 35
rect 1663 29 1673 31
rect 1675 35 1685 37
rect 1675 31 1679 35
rect 1683 31 1685 35
rect 1675 29 1685 31
rect 998 -101 1008 -99
rect 998 -105 1000 -101
rect 1004 -105 1008 -101
rect 998 -107 1008 -105
rect 1011 -107 1023 -99
rect 1026 -101 1036 -99
rect 1026 -105 1030 -101
rect 1034 -105 1036 -101
rect 1026 -107 1036 -105
rect 1066 -136 1076 -134
rect 931 -140 941 -138
rect 931 -144 933 -140
rect 937 -144 941 -140
rect 931 -146 941 -144
rect 944 -146 956 -138
rect 959 -140 969 -138
rect 959 -144 963 -140
rect 967 -144 969 -140
rect 1066 -140 1068 -136
rect 1072 -140 1076 -136
rect 1066 -142 1076 -140
rect 1079 -142 1091 -134
rect 1094 -136 1104 -134
rect 1094 -140 1098 -136
rect 1102 -140 1104 -136
rect 1094 -142 1104 -140
rect 959 -146 969 -144
rect 998 -184 1008 -182
rect 998 -188 1000 -184
rect 1004 -188 1008 -184
rect 998 -190 1008 -188
rect 1011 -190 1023 -182
rect 1026 -184 1036 -182
rect 1026 -188 1030 -184
rect 1034 -188 1036 -184
rect 1026 -190 1036 -188
rect 752 -285 762 -283
rect 752 -289 754 -285
rect 758 -289 762 -285
rect 752 -291 762 -289
rect 765 -291 777 -283
rect 780 -285 790 -283
rect 780 -289 784 -285
rect 788 -289 790 -285
rect 780 -291 790 -289
rect 987 -285 997 -283
rect 987 -289 989 -285
rect 993 -289 997 -285
rect 820 -320 830 -318
rect 685 -324 695 -322
rect 685 -328 687 -324
rect 691 -328 695 -324
rect 685 -330 695 -328
rect 698 -330 710 -322
rect 713 -324 723 -322
rect 713 -328 717 -324
rect 721 -328 723 -324
rect 820 -324 822 -320
rect 826 -324 830 -320
rect 820 -326 830 -324
rect 833 -326 845 -318
rect 848 -320 858 -318
rect 848 -324 852 -320
rect 856 -324 858 -320
rect 848 -326 858 -324
rect 713 -330 723 -328
rect 752 -368 762 -366
rect 752 -372 754 -368
rect 758 -372 762 -368
rect 752 -374 762 -372
rect 765 -374 777 -366
rect 780 -368 790 -366
rect 780 -372 784 -368
rect 788 -372 790 -368
rect 780 -374 790 -372
rect 666 -458 676 -456
rect 666 -462 668 -458
rect 672 -462 676 -458
rect 666 -464 676 -462
rect 679 -464 691 -456
rect 694 -458 704 -456
rect 694 -462 698 -458
rect 702 -462 704 -458
rect 694 -464 704 -462
rect 708 -458 718 -456
rect 708 -462 710 -458
rect 714 -462 718 -458
rect 708 -464 718 -462
rect 720 -458 730 -456
rect 720 -462 724 -458
rect 728 -462 730 -458
rect 720 -464 730 -462
rect 987 -291 997 -289
rect 1000 -291 1012 -283
rect 1015 -285 1025 -283
rect 1015 -289 1019 -285
rect 1023 -289 1025 -285
rect 1015 -291 1025 -289
rect 1055 -320 1065 -318
rect 920 -324 930 -322
rect 920 -328 922 -324
rect 926 -328 930 -324
rect 920 -330 930 -328
rect 933 -330 945 -322
rect 948 -324 958 -322
rect 948 -328 952 -324
rect 956 -328 958 -324
rect 1055 -324 1057 -320
rect 1061 -324 1065 -320
rect 1055 -326 1065 -324
rect 1068 -326 1080 -318
rect 1083 -320 1093 -318
rect 1083 -324 1087 -320
rect 1091 -324 1093 -320
rect 1083 -326 1093 -324
rect 948 -330 958 -328
rect 987 -368 997 -366
rect 987 -372 989 -368
rect 993 -372 997 -368
rect 987 -374 997 -372
rect 1000 -374 1012 -366
rect 1015 -368 1025 -366
rect 1015 -372 1019 -368
rect 1023 -372 1025 -368
rect 1015 -374 1025 -372
rect 918 -458 928 -456
rect 918 -462 920 -458
rect 924 -462 928 -458
rect 918 -464 928 -462
rect 931 -464 943 -456
rect 946 -458 956 -456
rect 946 -462 950 -458
rect 954 -462 956 -458
rect 946 -464 956 -462
rect 960 -458 970 -456
rect 960 -462 962 -458
rect 966 -462 970 -458
rect 960 -464 970 -462
rect 972 -458 982 -456
rect 972 -462 976 -458
rect 980 -462 982 -458
rect 972 -464 982 -462
rect 1035 -458 1045 -456
rect 1035 -462 1037 -458
rect 1041 -462 1045 -458
rect 1035 -464 1045 -462
rect 1048 -458 1060 -456
rect 1048 -462 1051 -458
rect 1055 -462 1060 -458
rect 1048 -464 1060 -462
rect 1063 -458 1073 -456
rect 1063 -462 1067 -458
rect 1071 -462 1073 -458
rect 1063 -464 1073 -462
rect 1077 -458 1087 -456
rect 1077 -462 1079 -458
rect 1083 -462 1087 -458
rect 1077 -464 1087 -462
rect 1089 -458 1099 -456
rect 1089 -462 1093 -458
rect 1097 -462 1099 -458
rect 1089 -464 1099 -462
rect 1975 35 1985 37
rect 1975 31 1977 35
rect 1981 31 1985 35
rect 1975 29 1985 31
rect 1988 29 2000 37
rect 2003 35 2013 37
rect 2003 31 2007 35
rect 2011 31 2013 35
rect 2003 29 2013 31
rect 2017 35 2027 37
rect 2017 31 2019 35
rect 2023 31 2027 35
rect 2017 29 2027 31
rect 2029 35 2039 37
rect 2029 31 2033 35
rect 2037 31 2039 35
rect 2029 29 2039 31
rect 2145 35 2155 37
rect 2145 31 2147 35
rect 2151 31 2155 35
rect 2145 29 2155 31
rect 2158 29 2170 37
rect 2173 35 2183 37
rect 2173 31 2177 35
rect 2181 31 2183 35
rect 2173 29 2183 31
rect 2187 35 2197 37
rect 2187 31 2189 35
rect 2193 31 2197 35
rect 2187 29 2197 31
rect 2199 35 2209 37
rect 2199 31 2203 35
rect 2207 31 2209 35
rect 2199 29 2209 31
rect 1504 -101 1514 -99
rect 1504 -105 1506 -101
rect 1510 -105 1514 -101
rect 1504 -107 1514 -105
rect 1517 -107 1529 -99
rect 1532 -101 1542 -99
rect 1532 -105 1536 -101
rect 1540 -105 1542 -101
rect 1532 -107 1542 -105
rect 1572 -136 1582 -134
rect 1437 -140 1447 -138
rect 1437 -144 1439 -140
rect 1443 -144 1447 -140
rect 1437 -146 1447 -144
rect 1450 -146 1462 -138
rect 1465 -140 1475 -138
rect 1465 -144 1469 -140
rect 1473 -144 1475 -140
rect 1572 -140 1574 -136
rect 1578 -140 1582 -136
rect 1572 -142 1582 -140
rect 1585 -142 1597 -134
rect 1600 -136 1610 -134
rect 1600 -140 1604 -136
rect 1608 -140 1610 -136
rect 1600 -142 1610 -140
rect 1465 -146 1475 -144
rect 1504 -184 1514 -182
rect 1504 -188 1506 -184
rect 1510 -188 1514 -184
rect 1504 -190 1514 -188
rect 1517 -190 1529 -182
rect 1532 -184 1542 -182
rect 1532 -188 1536 -184
rect 1540 -188 1542 -184
rect 1532 -190 1542 -188
rect 1275 -285 1285 -283
rect 1275 -289 1277 -285
rect 1281 -289 1285 -285
rect 1275 -291 1285 -289
rect 1288 -291 1300 -283
rect 1303 -285 1313 -283
rect 1303 -289 1307 -285
rect 1311 -289 1313 -285
rect 1303 -291 1313 -289
rect 1510 -285 1520 -283
rect 1510 -289 1512 -285
rect 1516 -289 1520 -285
rect 1343 -320 1353 -318
rect 1208 -324 1218 -322
rect 1208 -328 1210 -324
rect 1214 -328 1218 -324
rect 1208 -330 1218 -328
rect 1221 -330 1233 -322
rect 1236 -324 1246 -322
rect 1236 -328 1240 -324
rect 1244 -328 1246 -324
rect 1343 -324 1345 -320
rect 1349 -324 1353 -320
rect 1343 -326 1353 -324
rect 1356 -326 1368 -318
rect 1371 -320 1381 -318
rect 1371 -324 1375 -320
rect 1379 -324 1381 -320
rect 1371 -326 1381 -324
rect 1236 -330 1246 -328
rect 1275 -368 1285 -366
rect 1275 -372 1277 -368
rect 1281 -372 1285 -368
rect 1275 -374 1285 -372
rect 1288 -374 1300 -366
rect 1303 -368 1313 -366
rect 1303 -372 1307 -368
rect 1311 -372 1313 -368
rect 1303 -374 1313 -372
rect 1189 -458 1199 -456
rect 1189 -462 1191 -458
rect 1195 -462 1199 -458
rect 1189 -464 1199 -462
rect 1202 -464 1214 -456
rect 1217 -458 1227 -456
rect 1217 -462 1221 -458
rect 1225 -462 1227 -458
rect 1217 -464 1227 -462
rect 1231 -458 1241 -456
rect 1231 -462 1233 -458
rect 1237 -462 1241 -458
rect 1231 -464 1241 -462
rect 1243 -458 1253 -456
rect 1243 -462 1247 -458
rect 1251 -462 1253 -458
rect 1243 -464 1253 -462
rect 1510 -291 1520 -289
rect 1523 -291 1535 -283
rect 1538 -285 1548 -283
rect 1538 -289 1542 -285
rect 1546 -289 1548 -285
rect 1538 -291 1548 -289
rect 1578 -320 1588 -318
rect 1443 -324 1453 -322
rect 1443 -328 1445 -324
rect 1449 -328 1453 -324
rect 1443 -330 1453 -328
rect 1456 -330 1468 -322
rect 1471 -324 1481 -322
rect 1471 -328 1475 -324
rect 1479 -328 1481 -324
rect 1578 -324 1580 -320
rect 1584 -324 1588 -320
rect 1578 -326 1588 -324
rect 1591 -326 1603 -318
rect 1606 -320 1616 -318
rect 1606 -324 1610 -320
rect 1614 -324 1616 -320
rect 1606 -326 1616 -324
rect 1471 -330 1481 -328
rect 1510 -368 1520 -366
rect 1510 -372 1512 -368
rect 1516 -372 1520 -368
rect 1510 -374 1520 -372
rect 1523 -374 1535 -366
rect 1538 -368 1548 -366
rect 1538 -372 1542 -368
rect 1546 -372 1548 -368
rect 1538 -374 1548 -372
rect 1441 -458 1451 -456
rect 1441 -462 1443 -458
rect 1447 -462 1451 -458
rect 1441 -464 1451 -462
rect 1454 -464 1466 -456
rect 1469 -458 1479 -456
rect 1469 -462 1473 -458
rect 1477 -462 1479 -458
rect 1469 -464 1479 -462
rect 1483 -458 1493 -456
rect 1483 -462 1485 -458
rect 1489 -462 1493 -458
rect 1483 -464 1493 -462
rect 1495 -458 1505 -456
rect 1495 -462 1499 -458
rect 1503 -462 1505 -458
rect 1495 -464 1505 -462
rect 1558 -458 1568 -456
rect 1558 -462 1560 -458
rect 1564 -462 1568 -458
rect 1558 -464 1568 -462
rect 1571 -458 1583 -456
rect 1571 -462 1574 -458
rect 1578 -462 1583 -458
rect 1571 -464 1583 -462
rect 1586 -458 1596 -456
rect 1586 -462 1590 -458
rect 1594 -462 1596 -458
rect 1586 -464 1596 -462
rect 1600 -458 1610 -456
rect 1600 -462 1602 -458
rect 1606 -462 1610 -458
rect 1600 -464 1610 -462
rect 1612 -458 1622 -456
rect 1612 -462 1616 -458
rect 1620 -462 1622 -458
rect 1612 -464 1622 -462
rect 2028 -101 2038 -99
rect 2028 -105 2030 -101
rect 2034 -105 2038 -101
rect 2028 -107 2038 -105
rect 2041 -107 2053 -99
rect 2056 -101 2066 -99
rect 2056 -105 2060 -101
rect 2064 -105 2066 -101
rect 2056 -107 2066 -105
rect 2096 -136 2106 -134
rect 1961 -140 1971 -138
rect 1961 -144 1963 -140
rect 1967 -144 1971 -140
rect 1961 -146 1971 -144
rect 1974 -146 1986 -138
rect 1989 -140 1999 -138
rect 1989 -144 1993 -140
rect 1997 -144 1999 -140
rect 2096 -140 2098 -136
rect 2102 -140 2106 -136
rect 2096 -142 2106 -140
rect 2109 -142 2121 -134
rect 2124 -136 2134 -134
rect 2124 -140 2128 -136
rect 2132 -140 2134 -136
rect 2124 -142 2134 -140
rect 1989 -146 1999 -144
rect 2028 -184 2038 -182
rect 2028 -188 2030 -184
rect 2034 -188 2038 -184
rect 2028 -190 2038 -188
rect 2041 -190 2053 -182
rect 2056 -184 2066 -182
rect 2056 -188 2060 -184
rect 2064 -188 2066 -184
rect 2056 -190 2066 -188
rect 1798 -285 1808 -283
rect 1798 -289 1800 -285
rect 1804 -289 1808 -285
rect 1798 -291 1808 -289
rect 1811 -291 1823 -283
rect 1826 -285 1836 -283
rect 1826 -289 1830 -285
rect 1834 -289 1836 -285
rect 1826 -291 1836 -289
rect 2033 -285 2043 -283
rect 2033 -289 2035 -285
rect 2039 -289 2043 -285
rect 1866 -320 1876 -318
rect 1731 -324 1741 -322
rect 1731 -328 1733 -324
rect 1737 -328 1741 -324
rect 1731 -330 1741 -328
rect 1744 -330 1756 -322
rect 1759 -324 1769 -322
rect 1759 -328 1763 -324
rect 1767 -328 1769 -324
rect 1866 -324 1868 -320
rect 1872 -324 1876 -320
rect 1866 -326 1876 -324
rect 1879 -326 1891 -318
rect 1894 -320 1904 -318
rect 1894 -324 1898 -320
rect 1902 -324 1904 -320
rect 1894 -326 1904 -324
rect 1759 -330 1769 -328
rect 1798 -368 1808 -366
rect 1798 -372 1800 -368
rect 1804 -372 1808 -368
rect 1798 -374 1808 -372
rect 1811 -374 1823 -366
rect 1826 -368 1836 -366
rect 1826 -372 1830 -368
rect 1834 -372 1836 -368
rect 1826 -374 1836 -372
rect 1712 -458 1722 -456
rect 1712 -462 1714 -458
rect 1718 -462 1722 -458
rect 1712 -464 1722 -462
rect 1725 -464 1737 -456
rect 1740 -458 1750 -456
rect 1740 -462 1744 -458
rect 1748 -462 1750 -458
rect 1740 -464 1750 -462
rect 1754 -458 1764 -456
rect 1754 -462 1756 -458
rect 1760 -462 1764 -458
rect 1754 -464 1764 -462
rect 1766 -458 1776 -456
rect 1766 -462 1770 -458
rect 1774 -462 1776 -458
rect 1766 -464 1776 -462
rect 2033 -291 2043 -289
rect 2046 -291 2058 -283
rect 2061 -285 2071 -283
rect 2061 -289 2065 -285
rect 2069 -289 2071 -285
rect 2061 -291 2071 -289
rect 2101 -320 2111 -318
rect 1966 -324 1976 -322
rect 1966 -328 1968 -324
rect 1972 -328 1976 -324
rect 1966 -330 1976 -328
rect 1979 -330 1991 -322
rect 1994 -324 2004 -322
rect 1994 -328 1998 -324
rect 2002 -328 2004 -324
rect 2101 -324 2103 -320
rect 2107 -324 2111 -320
rect 2101 -326 2111 -324
rect 2114 -326 2126 -318
rect 2129 -320 2139 -318
rect 2129 -324 2133 -320
rect 2137 -324 2139 -320
rect 2129 -326 2139 -324
rect 1994 -330 2004 -328
rect 2033 -368 2043 -366
rect 2033 -372 2035 -368
rect 2039 -372 2043 -368
rect 2033 -374 2043 -372
rect 2046 -374 2058 -366
rect 2061 -368 2071 -366
rect 2061 -372 2065 -368
rect 2069 -372 2071 -368
rect 2061 -374 2071 -372
rect 1964 -458 1974 -456
rect 1964 -462 1966 -458
rect 1970 -462 1974 -458
rect 1964 -464 1974 -462
rect 1977 -464 1989 -456
rect 1992 -458 2002 -456
rect 1992 -462 1996 -458
rect 2000 -462 2002 -458
rect 1992 -464 2002 -462
rect 2006 -458 2016 -456
rect 2006 -462 2008 -458
rect 2012 -462 2016 -458
rect 2006 -464 2016 -462
rect 2018 -458 2028 -456
rect 2018 -462 2022 -458
rect 2026 -462 2028 -458
rect 2018 -464 2028 -462
rect 2081 -458 2091 -456
rect 2081 -462 2083 -458
rect 2087 -462 2091 -458
rect 2081 -464 2091 -462
rect 2094 -458 2106 -456
rect 2094 -462 2097 -458
rect 2101 -462 2106 -458
rect 2094 -464 2106 -462
rect 2109 -458 2119 -456
rect 2109 -462 2113 -458
rect 2117 -462 2119 -458
rect 2109 -464 2119 -462
rect 2123 -458 2133 -456
rect 2123 -462 2125 -458
rect 2129 -462 2133 -458
rect 2123 -464 2133 -462
rect 2135 -458 2145 -456
rect 2135 -462 2139 -458
rect 2143 -462 2145 -458
rect 2135 -464 2145 -462
rect 2321 -285 2331 -283
rect 2321 -289 2323 -285
rect 2327 -289 2331 -285
rect 2321 -291 2331 -289
rect 2334 -291 2346 -283
rect 2349 -285 2359 -283
rect 2349 -289 2353 -285
rect 2357 -289 2359 -285
rect 2349 -291 2359 -289
rect 2556 -285 2566 -283
rect 2556 -289 2558 -285
rect 2562 -289 2566 -285
rect 2389 -320 2399 -318
rect 2254 -324 2264 -322
rect 2254 -328 2256 -324
rect 2260 -328 2264 -324
rect 2254 -330 2264 -328
rect 2267 -330 2279 -322
rect 2282 -324 2292 -322
rect 2282 -328 2286 -324
rect 2290 -328 2292 -324
rect 2389 -324 2391 -320
rect 2395 -324 2399 -320
rect 2389 -326 2399 -324
rect 2402 -326 2414 -318
rect 2417 -320 2427 -318
rect 2417 -324 2421 -320
rect 2425 -324 2427 -320
rect 2417 -326 2427 -324
rect 2282 -330 2292 -328
rect 2321 -368 2331 -366
rect 2321 -372 2323 -368
rect 2327 -372 2331 -368
rect 2321 -374 2331 -372
rect 2334 -374 2346 -366
rect 2349 -368 2359 -366
rect 2349 -372 2353 -368
rect 2357 -372 2359 -368
rect 2349 -374 2359 -372
rect 2235 -458 2245 -456
rect 2235 -462 2237 -458
rect 2241 -462 2245 -458
rect 2235 -464 2245 -462
rect 2248 -464 2260 -456
rect 2263 -458 2273 -456
rect 2263 -462 2267 -458
rect 2271 -462 2273 -458
rect 2263 -464 2273 -462
rect 2277 -458 2287 -456
rect 2277 -462 2279 -458
rect 2283 -462 2287 -458
rect 2277 -464 2287 -462
rect 2289 -458 2299 -456
rect 2289 -462 2293 -458
rect 2297 -462 2299 -458
rect 2289 -464 2299 -462
rect 2556 -291 2566 -289
rect 2569 -291 2581 -283
rect 2584 -285 2594 -283
rect 2584 -289 2588 -285
rect 2592 -289 2594 -285
rect 2584 -291 2594 -289
rect 2624 -320 2634 -318
rect 2489 -324 2499 -322
rect 2489 -328 2491 -324
rect 2495 -328 2499 -324
rect 2489 -330 2499 -328
rect 2502 -330 2514 -322
rect 2517 -324 2527 -322
rect 2517 -328 2521 -324
rect 2525 -328 2527 -324
rect 2624 -324 2626 -320
rect 2630 -324 2634 -320
rect 2624 -326 2634 -324
rect 2637 -326 2649 -318
rect 2652 -320 2662 -318
rect 2652 -324 2656 -320
rect 2660 -324 2662 -320
rect 2652 -326 2662 -324
rect 2517 -330 2527 -328
rect 2556 -368 2566 -366
rect 2556 -372 2558 -368
rect 2562 -372 2566 -368
rect 2556 -374 2566 -372
rect 2569 -374 2581 -366
rect 2584 -368 2594 -366
rect 2584 -372 2588 -368
rect 2592 -372 2594 -368
rect 2584 -374 2594 -372
rect 2487 -458 2497 -456
rect 2487 -462 2489 -458
rect 2493 -462 2497 -458
rect 2487 -464 2497 -462
rect 2500 -464 2512 -456
rect 2515 -458 2525 -456
rect 2515 -462 2519 -458
rect 2523 -462 2525 -458
rect 2515 -464 2525 -462
rect 2529 -458 2539 -456
rect 2529 -462 2531 -458
rect 2535 -462 2539 -458
rect 2529 -464 2539 -462
rect 2541 -458 2551 -456
rect 2541 -462 2545 -458
rect 2549 -462 2551 -458
rect 2541 -464 2551 -462
rect 2604 -458 2614 -456
rect 2604 -462 2606 -458
rect 2610 -462 2614 -458
rect 2604 -464 2614 -462
rect 2617 -458 2629 -456
rect 2617 -462 2620 -458
rect 2624 -462 2629 -458
rect 2617 -464 2629 -462
rect 2632 -458 2642 -456
rect 2632 -462 2636 -458
rect 2640 -462 2642 -458
rect 2632 -464 2642 -462
rect 2646 -458 2656 -456
rect 2646 -462 2648 -458
rect 2652 -462 2656 -458
rect 2646 -464 2656 -462
rect 2658 -458 2668 -456
rect 2658 -462 2662 -458
rect 2666 -462 2668 -458
rect 2658 -464 2668 -462
<< pdiffusion >>
rect 8 1487 18 1489
rect 8 1483 10 1487
rect 14 1483 18 1487
rect 8 1481 18 1483
rect 20 1487 30 1489
rect 20 1483 24 1487
rect 28 1483 30 1487
rect 20 1481 30 1483
rect 34 1487 44 1489
rect 34 1483 36 1487
rect 40 1483 44 1487
rect 34 1481 44 1483
rect 47 1481 68 1489
rect 71 1481 94 1489
rect 97 1481 118 1489
rect 121 1487 131 1489
rect 121 1483 125 1487
rect 129 1483 131 1487
rect 121 1481 131 1483
rect 897 1303 907 1305
rect 897 1299 899 1303
rect 903 1299 907 1303
rect 897 1297 907 1299
rect 909 1303 919 1305
rect 909 1299 913 1303
rect 917 1299 919 1303
rect 909 1297 919 1299
rect 923 1303 933 1305
rect 923 1299 925 1303
rect 929 1299 933 1303
rect 923 1297 933 1299
rect 936 1303 948 1305
rect 936 1299 940 1303
rect 944 1299 948 1303
rect 936 1297 948 1299
rect 951 1303 961 1305
rect 951 1299 955 1303
rect 959 1299 961 1303
rect 951 1297 961 1299
rect 974 1303 984 1305
rect 974 1299 976 1303
rect 980 1299 984 1303
rect 974 1297 984 1299
rect 986 1303 996 1305
rect 986 1299 990 1303
rect 994 1299 996 1303
rect 986 1297 996 1299
rect 1000 1303 1010 1305
rect 1000 1299 1002 1303
rect 1006 1299 1010 1303
rect 1000 1297 1010 1299
rect 1013 1303 1025 1305
rect 1013 1299 1017 1303
rect 1021 1299 1025 1303
rect 1013 1297 1025 1299
rect 1028 1303 1038 1305
rect 1028 1299 1032 1303
rect 1036 1299 1038 1303
rect 1028 1297 1038 1299
rect 1042 1303 1052 1305
rect 1042 1299 1044 1303
rect 1048 1299 1052 1303
rect 1042 1297 1052 1299
rect 1054 1303 1064 1305
rect 1054 1299 1058 1303
rect 1062 1299 1064 1303
rect 1054 1297 1064 1299
rect 553 1288 563 1290
rect 196 1286 206 1288
rect 196 1282 198 1286
rect 202 1282 206 1286
rect 196 1280 206 1282
rect 208 1286 218 1288
rect 208 1282 212 1286
rect 216 1282 218 1286
rect 208 1280 218 1282
rect 222 1286 232 1288
rect 222 1282 224 1286
rect 228 1282 232 1286
rect 222 1280 232 1282
rect 235 1286 247 1288
rect 235 1282 239 1286
rect 243 1282 247 1286
rect 235 1280 247 1282
rect 250 1286 262 1288
rect 250 1282 254 1286
rect 258 1282 262 1286
rect 250 1280 262 1282
rect 265 1286 277 1288
rect 265 1282 269 1286
rect 273 1282 277 1286
rect 265 1280 277 1282
rect 280 1286 290 1288
rect 280 1282 284 1286
rect 288 1282 290 1286
rect 280 1280 290 1282
rect 303 1286 313 1288
rect 303 1282 305 1286
rect 309 1282 313 1286
rect 303 1280 313 1282
rect 315 1286 325 1288
rect 315 1282 319 1286
rect 323 1282 325 1286
rect 315 1280 325 1282
rect 329 1286 339 1288
rect 329 1282 331 1286
rect 335 1282 339 1286
rect 329 1280 339 1282
rect 342 1286 354 1288
rect 342 1282 346 1286
rect 350 1282 354 1286
rect 342 1280 354 1282
rect 357 1286 367 1288
rect 357 1282 361 1286
rect 365 1282 367 1286
rect 357 1280 367 1282
rect 371 1286 381 1288
rect 371 1282 373 1286
rect 377 1282 381 1286
rect 371 1280 381 1282
rect 383 1286 393 1288
rect 383 1282 387 1286
rect 391 1282 393 1286
rect 553 1284 555 1288
rect 559 1284 563 1288
rect 553 1282 563 1284
rect 565 1288 575 1290
rect 565 1284 569 1288
rect 573 1284 575 1288
rect 565 1282 575 1284
rect 579 1288 589 1290
rect 579 1284 581 1288
rect 585 1284 589 1288
rect 579 1282 589 1284
rect 592 1288 604 1290
rect 592 1284 596 1288
rect 600 1284 604 1288
rect 592 1282 604 1284
rect 607 1288 619 1290
rect 607 1284 611 1288
rect 615 1284 619 1288
rect 607 1282 619 1284
rect 622 1288 632 1290
rect 622 1284 626 1288
rect 630 1284 632 1288
rect 622 1282 632 1284
rect 649 1288 659 1290
rect 649 1284 651 1288
rect 655 1284 659 1288
rect 649 1282 659 1284
rect 661 1288 671 1290
rect 661 1284 665 1288
rect 669 1284 671 1288
rect 661 1282 671 1284
rect 675 1288 685 1290
rect 675 1284 677 1288
rect 681 1284 685 1288
rect 675 1282 685 1284
rect 688 1288 700 1290
rect 688 1284 692 1288
rect 696 1284 700 1288
rect 688 1282 700 1284
rect 703 1288 713 1290
rect 703 1284 707 1288
rect 711 1284 713 1288
rect 703 1282 713 1284
rect 717 1288 727 1290
rect 717 1284 719 1288
rect 723 1284 727 1288
rect 717 1282 727 1284
rect 729 1288 739 1290
rect 729 1284 733 1288
rect 737 1284 739 1288
rect 729 1282 739 1284
rect 383 1280 393 1282
rect 1304 1259 1314 1261
rect 1304 1255 1306 1259
rect 1310 1255 1314 1259
rect 1304 1253 1314 1255
rect 1316 1259 1326 1261
rect 1316 1255 1320 1259
rect 1324 1255 1326 1259
rect 1316 1253 1326 1255
rect 1330 1259 1340 1261
rect 1330 1255 1332 1259
rect 1336 1255 1340 1259
rect 1330 1253 1340 1255
rect 1343 1259 1355 1261
rect 1343 1255 1347 1259
rect 1351 1255 1355 1259
rect 1343 1253 1355 1255
rect 1358 1259 1368 1261
rect 1358 1255 1362 1259
rect 1366 1255 1368 1259
rect 1358 1253 1368 1255
rect 1372 1259 1382 1261
rect 1372 1255 1374 1259
rect 1378 1255 1382 1259
rect 1372 1253 1382 1255
rect 1384 1259 1394 1261
rect 1384 1255 1388 1259
rect 1392 1255 1394 1259
rect 1384 1253 1394 1255
rect 1334 1157 1344 1159
rect 988 1154 998 1156
rect 630 1149 640 1151
rect 630 1145 632 1149
rect 636 1145 640 1149
rect 286 1141 296 1143
rect 286 1137 288 1141
rect 292 1137 296 1141
rect 286 1135 296 1137
rect 299 1141 311 1143
rect 299 1137 303 1141
rect 307 1137 311 1141
rect 299 1135 311 1137
rect 314 1141 324 1143
rect 314 1137 318 1141
rect 322 1137 324 1141
rect 630 1143 640 1145
rect 643 1149 655 1151
rect 643 1145 647 1149
rect 651 1145 655 1149
rect 643 1143 655 1145
rect 658 1149 668 1151
rect 988 1150 990 1154
rect 994 1150 998 1154
rect 658 1145 662 1149
rect 666 1145 668 1149
rect 658 1143 668 1145
rect 314 1135 324 1137
rect 988 1148 998 1150
rect 1001 1154 1013 1156
rect 1001 1150 1005 1154
rect 1009 1150 1013 1154
rect 1001 1148 1013 1150
rect 1016 1154 1026 1156
rect 1016 1150 1020 1154
rect 1024 1150 1026 1154
rect 1334 1153 1336 1157
rect 1340 1153 1344 1157
rect 1016 1148 1026 1150
rect 1334 1151 1344 1153
rect 1347 1157 1359 1159
rect 1347 1153 1351 1157
rect 1355 1153 1359 1157
rect 1347 1151 1359 1153
rect 1362 1157 1372 1159
rect 1362 1153 1366 1157
rect 1370 1153 1372 1157
rect 1362 1151 1372 1153
rect 161 1102 171 1104
rect 161 1098 163 1102
rect 167 1098 171 1102
rect 161 1096 171 1098
rect 173 1102 183 1104
rect 173 1098 177 1102
rect 181 1098 183 1102
rect 173 1096 183 1098
rect 218 1093 228 1095
rect 218 1089 220 1093
rect 224 1089 228 1093
rect 218 1087 228 1089
rect 231 1093 243 1095
rect 231 1089 235 1093
rect 239 1089 243 1093
rect 231 1087 243 1089
rect 246 1093 256 1095
rect 246 1089 250 1093
rect 254 1089 256 1093
rect 505 1110 515 1112
rect 505 1106 507 1110
rect 511 1106 515 1110
rect 505 1104 515 1106
rect 517 1110 527 1112
rect 517 1106 521 1110
rect 525 1106 527 1110
rect 517 1104 527 1106
rect 562 1101 572 1103
rect 353 1097 363 1099
rect 353 1093 355 1097
rect 359 1093 363 1097
rect 246 1087 256 1089
rect 353 1091 363 1093
rect 366 1097 378 1099
rect 366 1093 370 1097
rect 374 1093 378 1097
rect 366 1091 378 1093
rect 381 1097 391 1099
rect 381 1093 385 1097
rect 389 1093 391 1097
rect 562 1097 564 1101
rect 568 1097 572 1101
rect 381 1091 391 1093
rect 562 1095 572 1097
rect 575 1101 587 1103
rect 575 1097 579 1101
rect 583 1097 587 1101
rect 575 1095 587 1097
rect 590 1101 600 1103
rect 590 1097 594 1101
rect 598 1097 600 1101
rect 863 1115 873 1117
rect 863 1111 865 1115
rect 869 1111 873 1115
rect 863 1109 873 1111
rect 875 1115 885 1117
rect 875 1111 879 1115
rect 883 1111 885 1115
rect 875 1109 885 1111
rect 697 1105 707 1107
rect 697 1101 699 1105
rect 703 1101 707 1105
rect 590 1095 600 1097
rect 697 1099 707 1101
rect 710 1105 722 1107
rect 710 1101 714 1105
rect 718 1101 722 1105
rect 710 1099 722 1101
rect 725 1105 735 1107
rect 920 1106 930 1108
rect 725 1101 729 1105
rect 733 1101 735 1105
rect 920 1102 922 1106
rect 926 1102 930 1106
rect 725 1099 735 1101
rect 920 1100 930 1102
rect 933 1106 945 1108
rect 933 1102 937 1106
rect 941 1102 945 1106
rect 933 1100 945 1102
rect 948 1106 958 1108
rect 948 1102 952 1106
rect 956 1102 958 1106
rect 1209 1118 1219 1120
rect 1209 1114 1211 1118
rect 1215 1114 1219 1118
rect 1209 1112 1219 1114
rect 1221 1118 1231 1120
rect 1221 1114 1225 1118
rect 1229 1114 1231 1118
rect 1221 1112 1231 1114
rect 1055 1110 1065 1112
rect 1055 1106 1057 1110
rect 1061 1106 1065 1110
rect 948 1100 958 1102
rect 1055 1104 1065 1106
rect 1068 1110 1080 1112
rect 1068 1106 1072 1110
rect 1076 1106 1080 1110
rect 1068 1104 1080 1106
rect 1083 1110 1093 1112
rect 1083 1106 1087 1110
rect 1091 1106 1093 1110
rect 1266 1109 1276 1111
rect 1083 1104 1093 1106
rect 1266 1105 1268 1109
rect 1272 1105 1276 1109
rect 1266 1103 1276 1105
rect 1279 1109 1291 1111
rect 1279 1105 1283 1109
rect 1287 1105 1291 1109
rect 1279 1103 1291 1105
rect 1294 1109 1304 1111
rect 1294 1105 1298 1109
rect 1302 1105 1304 1109
rect 1401 1113 1411 1115
rect 1401 1109 1403 1113
rect 1407 1109 1411 1113
rect 1294 1103 1304 1105
rect 1401 1107 1411 1109
rect 1414 1113 1426 1115
rect 1414 1109 1418 1113
rect 1422 1109 1426 1113
rect 1414 1107 1426 1109
rect 1429 1113 1439 1115
rect 1429 1109 1433 1113
rect 1437 1109 1439 1113
rect 1429 1107 1439 1109
rect 1334 1074 1344 1076
rect 988 1071 998 1073
rect 630 1066 640 1068
rect 630 1062 632 1066
rect 636 1062 640 1066
rect 630 1060 640 1062
rect 643 1066 655 1068
rect 643 1062 647 1066
rect 651 1062 655 1066
rect 643 1060 655 1062
rect 658 1066 668 1068
rect 658 1062 662 1066
rect 666 1062 668 1066
rect 988 1067 990 1071
rect 994 1067 998 1071
rect 988 1065 998 1067
rect 1001 1071 1013 1073
rect 1001 1067 1005 1071
rect 1009 1067 1013 1071
rect 1001 1065 1013 1067
rect 1016 1071 1026 1073
rect 1016 1067 1020 1071
rect 1024 1067 1026 1071
rect 1334 1070 1336 1074
rect 1340 1070 1344 1074
rect 1334 1068 1344 1070
rect 1347 1074 1359 1076
rect 1347 1070 1351 1074
rect 1355 1070 1359 1074
rect 1347 1068 1359 1070
rect 1362 1074 1372 1076
rect 1362 1070 1366 1074
rect 1370 1070 1372 1074
rect 1362 1068 1372 1070
rect 1016 1065 1026 1067
rect 658 1060 668 1062
rect 286 1058 296 1060
rect 286 1054 288 1058
rect 292 1054 296 1058
rect 286 1052 296 1054
rect 299 1058 311 1060
rect 299 1054 303 1058
rect 307 1054 311 1058
rect 299 1052 311 1054
rect 314 1058 324 1060
rect 314 1054 318 1058
rect 322 1054 324 1058
rect 314 1052 324 1054
rect -97 988 -87 990
rect -97 984 -95 988
rect -91 984 -87 988
rect -97 982 -87 984
rect -85 988 -75 990
rect -85 984 -81 988
rect -77 984 -75 988
rect -85 982 -75 984
rect -71 988 -61 990
rect -71 984 -69 988
rect -65 984 -61 988
rect -71 982 -61 984
rect -58 988 -46 990
rect -58 984 -54 988
rect -50 984 -46 988
rect -58 982 -46 984
rect -43 988 -31 990
rect -43 984 -39 988
rect -35 984 -31 988
rect -43 982 -31 984
rect -28 988 -16 990
rect -28 984 -24 988
rect -20 984 -16 988
rect -28 982 -16 984
rect -13 988 -3 990
rect -13 984 -9 988
rect -5 984 -3 988
rect -13 982 -3 984
rect 1312 979 1322 981
rect 1312 975 1314 979
rect 1318 975 1322 979
rect 1312 973 1322 975
rect 1324 979 1334 981
rect 1324 975 1328 979
rect 1332 975 1334 979
rect 1324 973 1334 975
rect 1338 979 1348 981
rect 1338 975 1340 979
rect 1344 975 1348 979
rect 1338 973 1348 975
rect 1351 979 1363 981
rect 1351 975 1355 979
rect 1359 975 1363 979
rect 1351 973 1363 975
rect 1366 979 1376 981
rect 1366 975 1370 979
rect 1374 975 1376 979
rect 1366 973 1376 975
rect 1380 979 1390 981
rect 1380 975 1382 979
rect 1386 975 1390 979
rect 1380 973 1390 975
rect 1392 979 1402 981
rect 1392 975 1396 979
rect 1400 975 1402 979
rect 1392 973 1402 975
rect 889 936 899 938
rect 889 932 891 936
rect 895 932 899 936
rect 889 930 899 932
rect 901 936 911 938
rect 901 932 905 936
rect 909 932 911 936
rect 901 930 911 932
rect 915 936 925 938
rect 915 932 917 936
rect 921 932 925 936
rect 915 930 925 932
rect 928 936 940 938
rect 928 932 932 936
rect 936 932 940 936
rect 928 930 940 932
rect 943 936 953 938
rect 943 932 947 936
rect 951 932 953 936
rect 943 930 953 932
rect 966 936 976 938
rect 966 932 968 936
rect 972 932 976 936
rect 966 930 976 932
rect 978 936 988 938
rect 978 932 982 936
rect 986 932 988 936
rect 978 930 988 932
rect 992 936 1002 938
rect 992 932 994 936
rect 998 932 1002 936
rect 992 930 1002 932
rect 1005 936 1017 938
rect 1005 932 1009 936
rect 1013 932 1017 936
rect 1005 930 1017 932
rect 1020 936 1030 938
rect 1020 932 1024 936
rect 1028 932 1030 936
rect 1020 930 1030 932
rect 1034 936 1044 938
rect 1034 932 1036 936
rect 1040 932 1044 936
rect 1034 930 1044 932
rect 1046 936 1056 938
rect 1046 932 1050 936
rect 1054 932 1056 936
rect 1046 930 1056 932
rect 525 923 535 925
rect 525 919 527 923
rect 531 919 535 923
rect 525 917 535 919
rect 537 923 547 925
rect 537 919 541 923
rect 545 919 547 923
rect 537 917 547 919
rect 551 923 561 925
rect 551 919 553 923
rect 557 919 561 923
rect 551 917 561 919
rect 564 923 576 925
rect 564 919 568 923
rect 572 919 576 923
rect 564 917 576 919
rect 579 923 591 925
rect 579 919 583 923
rect 587 919 591 923
rect 579 917 591 919
rect 594 923 604 925
rect 594 919 598 923
rect 602 919 604 923
rect 594 917 604 919
rect 621 923 631 925
rect 621 919 623 923
rect 627 919 631 923
rect 621 917 631 919
rect 633 923 643 925
rect 633 919 637 923
rect 641 919 643 923
rect 633 917 643 919
rect 647 923 657 925
rect 647 919 649 923
rect 653 919 657 923
rect 647 917 657 919
rect 660 923 672 925
rect 660 919 664 923
rect 668 919 672 923
rect 660 917 672 919
rect 675 923 685 925
rect 675 919 679 923
rect 683 919 685 923
rect 675 917 685 919
rect 689 923 699 925
rect 689 919 691 923
rect 695 919 699 923
rect 689 917 699 919
rect 701 923 711 925
rect 701 919 705 923
rect 709 919 711 923
rect 701 917 711 919
rect 182 915 192 917
rect 182 911 184 915
rect 188 911 192 915
rect 182 909 192 911
rect 194 915 204 917
rect 194 911 198 915
rect 202 911 204 915
rect 194 909 204 911
rect 208 915 218 917
rect 208 911 210 915
rect 214 911 218 915
rect 208 909 218 911
rect 221 915 233 917
rect 221 911 225 915
rect 229 911 233 915
rect 221 909 233 911
rect 236 915 248 917
rect 236 911 240 915
rect 244 911 248 915
rect 236 909 248 911
rect 251 915 263 917
rect 251 911 255 915
rect 259 911 263 915
rect 251 909 263 911
rect 266 915 276 917
rect 266 911 270 915
rect 274 911 276 915
rect 266 909 276 911
rect 289 915 299 917
rect 289 911 291 915
rect 295 911 299 915
rect 289 909 299 911
rect 301 915 311 917
rect 301 911 305 915
rect 309 911 311 915
rect 301 909 311 911
rect 315 915 325 917
rect 315 911 317 915
rect 321 911 325 915
rect 315 909 325 911
rect 328 915 340 917
rect 328 911 332 915
rect 336 911 340 915
rect 328 909 340 911
rect 343 915 353 917
rect 343 911 347 915
rect 351 911 353 915
rect 343 909 353 911
rect 357 915 367 917
rect 357 911 359 915
rect 363 911 367 915
rect 357 909 367 911
rect 369 915 379 917
rect 369 911 373 915
rect 377 911 379 915
rect 369 909 379 911
rect -45 824 -35 826
rect -45 820 -43 824
rect -39 820 -35 824
rect -45 818 -35 820
rect -33 824 -23 826
rect -33 820 -29 824
rect -25 820 -23 824
rect -33 818 -23 820
rect -19 824 -9 826
rect -19 820 -17 824
rect -13 820 -9 824
rect -19 818 -9 820
rect -6 818 15 826
rect 18 818 41 826
rect 44 818 65 826
rect 68 824 78 826
rect 68 820 72 824
rect 76 820 78 824
rect 68 818 78 820
rect 133 265 143 267
rect 133 261 135 265
rect 139 261 143 265
rect 133 259 143 261
rect 146 265 158 267
rect 146 261 150 265
rect 154 261 158 265
rect 146 259 158 261
rect 161 265 171 267
rect 161 261 165 265
rect 169 261 171 265
rect 161 259 171 261
rect 175 265 185 267
rect 175 261 177 265
rect 181 261 185 265
rect 175 259 185 261
rect 187 265 197 267
rect 187 261 191 265
rect 195 261 197 265
rect 187 259 197 261
rect -794 204 -784 206
rect -794 200 -792 204
rect -788 200 -784 204
rect -794 198 -784 200
rect -781 204 -769 206
rect -781 200 -777 204
rect -773 200 -769 204
rect -781 198 -769 200
rect -766 204 -756 206
rect -766 200 -762 204
rect -758 200 -756 204
rect -766 198 -756 200
rect -752 204 -742 206
rect -752 200 -750 204
rect -746 200 -742 204
rect -752 198 -742 200
rect -740 204 -730 206
rect -740 200 -736 204
rect -732 200 -730 204
rect -740 198 -730 200
rect -717 204 -707 206
rect -717 200 -715 204
rect -711 200 -707 204
rect -717 198 -707 200
rect -704 204 -692 206
rect -704 200 -700 204
rect -696 200 -692 204
rect -704 198 -692 200
rect -689 204 -679 206
rect -689 200 -685 204
rect -681 200 -679 204
rect -689 198 -679 200
rect -675 204 -665 206
rect -675 200 -673 204
rect -669 200 -665 204
rect -675 198 -665 200
rect -663 204 -653 206
rect -663 200 -659 204
rect -655 200 -653 204
rect -663 198 -653 200
rect -640 204 -630 206
rect -640 200 -638 204
rect -634 200 -630 204
rect -640 198 -630 200
rect -627 204 -615 206
rect -627 200 -623 204
rect -619 200 -615 204
rect -627 198 -615 200
rect -612 204 -602 206
rect -612 200 -608 204
rect -604 200 -602 204
rect -612 198 -602 200
rect -598 204 -588 206
rect -598 200 -596 204
rect -592 200 -588 204
rect -598 198 -588 200
rect -586 204 -576 206
rect -586 200 -582 204
rect -578 200 -576 204
rect -586 198 -576 200
rect -563 204 -553 206
rect -563 200 -561 204
rect -557 200 -553 204
rect -563 198 -553 200
rect -550 204 -538 206
rect -550 200 -546 204
rect -542 200 -538 204
rect -550 198 -538 200
rect -535 204 -525 206
rect -535 200 -531 204
rect -527 200 -525 204
rect -535 198 -525 200
rect -521 204 -511 206
rect -521 200 -519 204
rect -515 200 -511 204
rect -521 198 -511 200
rect -509 204 -499 206
rect -509 200 -505 204
rect -501 200 -499 204
rect -509 198 -499 200
rect -486 204 -476 206
rect -486 200 -484 204
rect -480 200 -476 204
rect -486 198 -476 200
rect -473 204 -461 206
rect -473 200 -469 204
rect -465 200 -461 204
rect -473 198 -461 200
rect -458 204 -448 206
rect -458 200 -454 204
rect -450 200 -448 204
rect -458 198 -448 200
rect -444 204 -434 206
rect -444 200 -442 204
rect -438 200 -434 204
rect -444 198 -434 200
rect -432 204 -422 206
rect -432 200 -428 204
rect -424 200 -422 204
rect -432 198 -422 200
rect -409 204 -399 206
rect -409 200 -407 204
rect -403 200 -399 204
rect -409 198 -399 200
rect -396 204 -384 206
rect -396 200 -392 204
rect -388 200 -384 204
rect -396 198 -384 200
rect -381 204 -371 206
rect -381 200 -377 204
rect -373 200 -371 204
rect -381 198 -371 200
rect -367 204 -357 206
rect -367 200 -365 204
rect -361 200 -357 204
rect -367 198 -357 200
rect -355 204 -345 206
rect -355 200 -351 204
rect -347 200 -345 204
rect -355 198 -345 200
rect -332 204 -322 206
rect -332 200 -330 204
rect -326 200 -322 204
rect -332 198 -322 200
rect -319 204 -307 206
rect -319 200 -315 204
rect -311 200 -307 204
rect -319 198 -307 200
rect -304 204 -294 206
rect -304 200 -300 204
rect -296 200 -294 204
rect -304 198 -294 200
rect -290 204 -280 206
rect -290 200 -288 204
rect -284 200 -280 204
rect -290 198 -280 200
rect -278 204 -268 206
rect -278 200 -274 204
rect -270 200 -268 204
rect -278 198 -268 200
rect -255 204 -245 206
rect -255 200 -253 204
rect -249 200 -245 204
rect -255 198 -245 200
rect -242 204 -230 206
rect -242 200 -238 204
rect -234 200 -230 204
rect -242 198 -230 200
rect -227 204 -217 206
rect -227 200 -223 204
rect -219 200 -217 204
rect -227 198 -217 200
rect -213 204 -203 206
rect -213 200 -211 204
rect -207 200 -203 204
rect -213 198 -203 200
rect -201 204 -191 206
rect -201 200 -197 204
rect -193 200 -191 204
rect -201 198 -191 200
rect -73 189 -63 191
rect -73 185 -71 189
rect -67 185 -63 189
rect -73 183 -63 185
rect -61 189 -51 191
rect -61 185 -57 189
rect -53 185 -51 189
rect -61 183 -51 185
rect -73 105 -63 107
rect -73 101 -71 105
rect -67 101 -63 105
rect -73 99 -63 101
rect -61 105 -51 107
rect -61 101 -57 105
rect -53 101 -51 105
rect -61 99 -51 101
rect 135 189 145 191
rect 135 185 137 189
rect 141 185 145 189
rect 135 183 145 185
rect 148 189 160 191
rect 148 185 152 189
rect 156 185 160 189
rect 148 183 160 185
rect 163 189 173 191
rect 163 185 167 189
rect 171 185 173 189
rect 163 183 173 185
rect 177 189 187 191
rect 177 185 179 189
rect 183 185 187 189
rect 177 183 187 185
rect 189 189 199 191
rect 189 185 193 189
rect 197 185 199 189
rect 189 183 199 185
rect 281 189 291 191
rect 281 185 283 189
rect 287 185 291 189
rect 281 183 291 185
rect 294 189 306 191
rect 294 185 298 189
rect 302 185 306 189
rect 294 183 306 185
rect 309 189 319 191
rect 309 185 313 189
rect 317 185 319 189
rect 309 183 319 185
rect 323 189 333 191
rect 323 185 325 189
rect 329 185 333 189
rect 323 183 333 185
rect 335 189 345 191
rect 335 185 339 189
rect 343 185 345 189
rect 335 183 345 185
rect 451 189 461 191
rect 451 185 453 189
rect 457 185 461 189
rect 451 183 461 185
rect 464 189 476 191
rect 464 185 468 189
rect 472 185 476 189
rect 464 183 476 185
rect 479 189 489 191
rect 479 185 483 189
rect 487 185 489 189
rect 479 183 489 185
rect 493 189 503 191
rect 493 185 495 189
rect 499 185 503 189
rect 493 183 503 185
rect 505 189 515 191
rect 505 185 509 189
rect 513 185 515 189
rect 505 183 515 185
rect 839 189 849 191
rect 839 185 841 189
rect 845 185 849 189
rect 839 183 849 185
rect 852 189 864 191
rect 852 185 856 189
rect 860 185 864 189
rect 852 183 864 185
rect 867 189 877 191
rect 867 185 871 189
rect 875 185 877 189
rect 867 183 877 185
rect 881 189 891 191
rect 881 185 883 189
rect 887 185 891 189
rect 881 183 891 185
rect 893 189 903 191
rect 893 185 897 189
rect 901 185 903 189
rect 893 183 903 185
rect 1009 189 1019 191
rect 1009 185 1011 189
rect 1015 185 1019 189
rect 1009 183 1019 185
rect 1022 189 1034 191
rect 1022 185 1026 189
rect 1030 185 1034 189
rect 1022 183 1034 185
rect 1037 189 1047 191
rect 1037 185 1041 189
rect 1045 185 1047 189
rect 1037 183 1047 185
rect 1051 189 1061 191
rect 1051 185 1053 189
rect 1057 185 1061 189
rect 1051 183 1061 185
rect 1063 189 1073 191
rect 1063 185 1067 189
rect 1071 185 1073 189
rect 1063 183 1073 185
rect 1344 189 1354 191
rect 1344 185 1346 189
rect 1350 185 1354 189
rect 1344 183 1354 185
rect 1357 189 1369 191
rect 1357 185 1361 189
rect 1365 185 1369 189
rect 1357 183 1369 185
rect 1372 189 1382 191
rect 1372 185 1376 189
rect 1380 185 1382 189
rect 1372 183 1382 185
rect 1386 189 1396 191
rect 1386 185 1388 189
rect 1392 185 1396 189
rect 1386 183 1396 185
rect 1398 189 1408 191
rect 1398 185 1402 189
rect 1406 185 1408 189
rect 1398 183 1408 185
rect 1514 189 1524 191
rect 1514 185 1516 189
rect 1520 185 1524 189
rect 1514 183 1524 185
rect 1527 189 1539 191
rect 1527 185 1531 189
rect 1535 185 1539 189
rect 1527 183 1539 185
rect 1542 189 1552 191
rect 1542 185 1546 189
rect 1550 185 1552 189
rect 1542 183 1552 185
rect 1556 189 1566 191
rect 1556 185 1558 189
rect 1562 185 1566 189
rect 1556 183 1566 185
rect 1568 189 1578 191
rect 1568 185 1572 189
rect 1576 185 1578 189
rect 1568 183 1578 185
rect 1868 189 1878 191
rect 1868 185 1870 189
rect 1874 185 1878 189
rect 1868 183 1878 185
rect 1881 189 1893 191
rect 1881 185 1885 189
rect 1889 185 1893 189
rect 1881 183 1893 185
rect 1896 189 1906 191
rect 1896 185 1900 189
rect 1904 185 1906 189
rect 1896 183 1906 185
rect 1910 189 1920 191
rect 1910 185 1912 189
rect 1916 185 1920 189
rect 1910 183 1920 185
rect 1922 189 1932 191
rect 1922 185 1926 189
rect 1930 185 1932 189
rect 1922 183 1932 185
rect 2038 189 2048 191
rect 2038 185 2040 189
rect 2044 185 2048 189
rect 2038 183 2048 185
rect 2051 189 2063 191
rect 2051 185 2055 189
rect 2059 185 2063 189
rect 2051 183 2063 185
rect 2066 189 2076 191
rect 2066 185 2070 189
rect 2074 185 2076 189
rect 2066 183 2076 185
rect 2080 189 2090 191
rect 2080 185 2082 189
rect 2086 185 2090 189
rect 2080 183 2090 185
rect 2092 189 2102 191
rect 2092 185 2096 189
rect 2100 185 2102 189
rect 2092 183 2102 185
rect 137 113 147 115
rect 137 109 139 113
rect 143 109 147 113
rect 137 107 147 109
rect 150 113 162 115
rect 150 109 154 113
rect 158 109 162 113
rect 150 107 162 109
rect 165 113 175 115
rect 165 109 169 113
rect 173 109 175 113
rect 165 107 175 109
rect 179 113 189 115
rect 179 109 181 113
rect 185 109 189 113
rect 179 107 189 109
rect 191 113 201 115
rect 191 109 195 113
rect 199 109 201 113
rect 191 107 201 109
rect -619 25 -609 27
rect -619 21 -617 25
rect -613 21 -609 25
rect -619 19 -609 21
rect -606 25 -594 27
rect -606 21 -602 25
rect -598 21 -594 25
rect -606 19 -594 21
rect -591 25 -581 27
rect -591 21 -587 25
rect -583 21 -581 25
rect -591 19 -581 21
rect -577 25 -567 27
rect -577 21 -575 25
rect -571 21 -567 25
rect -577 19 -567 21
rect -565 25 -555 27
rect -565 21 -561 25
rect -557 21 -555 25
rect -565 19 -555 21
rect -542 25 -532 27
rect -542 21 -540 25
rect -536 21 -532 25
rect -542 19 -532 21
rect -529 25 -517 27
rect -529 21 -525 25
rect -521 21 -517 25
rect -529 19 -517 21
rect -514 25 -504 27
rect -514 21 -510 25
rect -506 21 -504 25
rect -514 19 -504 21
rect -500 25 -490 27
rect -500 21 -498 25
rect -494 21 -490 25
rect -500 19 -490 21
rect -488 25 -478 27
rect -488 21 -484 25
rect -480 21 -478 25
rect -488 19 -478 21
rect -465 25 -455 27
rect -465 21 -463 25
rect -459 21 -455 25
rect -465 19 -455 21
rect -452 25 -440 27
rect -452 21 -448 25
rect -444 21 -440 25
rect -452 19 -440 21
rect -437 25 -427 27
rect -437 21 -433 25
rect -429 21 -427 25
rect -437 19 -427 21
rect -423 25 -413 27
rect -423 21 -421 25
rect -417 21 -413 25
rect -423 19 -413 21
rect -411 25 -401 27
rect -411 21 -407 25
rect -403 21 -401 25
rect -411 19 -401 21
rect -388 25 -378 27
rect -388 21 -386 25
rect -382 21 -378 25
rect -388 19 -378 21
rect -375 25 -363 27
rect -375 21 -371 25
rect -367 21 -363 25
rect -375 19 -363 21
rect -360 25 -350 27
rect -360 21 -356 25
rect -352 21 -350 25
rect -360 19 -350 21
rect -346 25 -336 27
rect -346 21 -344 25
rect -340 21 -336 25
rect -346 19 -336 21
rect -334 25 -324 27
rect -334 21 -330 25
rect -326 21 -324 25
rect -334 19 -324 21
rect 266 75 276 77
rect 266 71 268 75
rect 272 71 276 75
rect 266 69 276 71
rect 279 69 291 77
rect 294 75 304 77
rect 294 71 298 75
rect 302 71 304 75
rect 294 69 304 71
rect 308 75 318 77
rect 308 71 310 75
rect 314 71 318 75
rect 308 69 318 71
rect 320 75 330 77
rect 320 71 324 75
rect 328 71 330 75
rect 320 69 330 71
rect 139 37 149 39
rect 139 33 141 37
rect 145 33 149 37
rect 139 31 149 33
rect 152 37 164 39
rect 152 33 156 37
rect 160 33 164 37
rect 152 31 164 33
rect 167 37 177 39
rect 167 33 171 37
rect 175 33 177 37
rect 167 31 177 33
rect 181 37 191 39
rect 181 33 183 37
rect 187 33 191 37
rect 181 31 191 33
rect 193 37 203 39
rect 388 75 398 77
rect 388 71 390 75
rect 394 71 398 75
rect 388 69 398 71
rect 401 75 413 77
rect 401 71 405 75
rect 409 71 413 75
rect 401 69 413 71
rect 416 75 426 77
rect 416 71 420 75
rect 424 71 426 75
rect 416 69 426 71
rect 430 75 440 77
rect 430 71 432 75
rect 436 71 440 75
rect 430 69 440 71
rect 442 75 452 77
rect 442 71 446 75
rect 450 71 452 75
rect 442 69 452 71
rect 558 75 568 77
rect 558 71 560 75
rect 564 71 568 75
rect 558 69 568 71
rect 571 75 583 77
rect 571 71 575 75
rect 579 71 583 75
rect 571 69 583 71
rect 586 75 596 77
rect 586 71 590 75
rect 594 71 596 75
rect 586 69 596 71
rect 600 75 610 77
rect 600 71 602 75
rect 606 71 610 75
rect 600 69 610 71
rect 612 75 622 77
rect 612 71 616 75
rect 620 71 622 75
rect 612 69 622 71
rect 193 33 197 37
rect 201 33 203 37
rect 193 31 203 33
rect 946 75 956 77
rect 946 71 948 75
rect 952 71 956 75
rect 946 69 956 71
rect 959 75 971 77
rect 959 71 963 75
rect 967 71 971 75
rect 959 69 971 71
rect 974 75 984 77
rect 974 71 978 75
rect 982 71 984 75
rect 974 69 984 71
rect 988 75 998 77
rect 988 71 990 75
rect 994 71 998 75
rect 988 69 998 71
rect 1000 75 1010 77
rect 1000 71 1004 75
rect 1008 71 1010 75
rect 1000 69 1010 71
rect 485 -61 495 -59
rect 485 -65 487 -61
rect 491 -65 495 -61
rect 485 -67 495 -65
rect 498 -61 510 -59
rect 498 -65 502 -61
rect 506 -65 510 -61
rect 498 -67 510 -65
rect 513 -61 523 -59
rect 513 -65 517 -61
rect 521 -65 523 -61
rect 513 -67 523 -65
rect 418 -100 428 -98
rect 418 -104 420 -100
rect 424 -104 428 -100
rect 418 -106 428 -104
rect 431 -100 443 -98
rect 431 -104 435 -100
rect 439 -104 443 -100
rect 431 -106 443 -104
rect 446 -100 456 -98
rect 553 -96 563 -94
rect 446 -104 450 -100
rect 454 -104 456 -100
rect 446 -106 456 -104
rect 553 -100 555 -96
rect 559 -100 563 -96
rect 553 -102 563 -100
rect 566 -96 578 -94
rect 566 -100 570 -96
rect 574 -100 578 -96
rect 566 -102 578 -100
rect 581 -96 591 -94
rect 581 -100 585 -96
rect 589 -100 591 -96
rect 581 -102 591 -100
rect 485 -144 495 -142
rect 485 -148 487 -144
rect 491 -148 495 -144
rect 485 -150 495 -148
rect 498 -144 510 -142
rect 498 -148 502 -144
rect 506 -148 510 -144
rect 498 -150 510 -148
rect 513 -144 523 -142
rect 513 -148 517 -144
rect 521 -148 523 -144
rect 513 -150 523 -148
rect 1116 75 1126 77
rect 1116 71 1118 75
rect 1122 71 1126 75
rect 1116 69 1126 71
rect 1129 75 1141 77
rect 1129 71 1133 75
rect 1137 71 1141 75
rect 1129 69 1141 71
rect 1144 75 1154 77
rect 1144 71 1148 75
rect 1152 71 1154 75
rect 1144 69 1154 71
rect 1158 75 1168 77
rect 1158 71 1160 75
rect 1164 71 1168 75
rect 1158 69 1168 71
rect 1170 75 1180 77
rect 1170 71 1174 75
rect 1178 71 1180 75
rect 1170 69 1180 71
rect 1451 75 1461 77
rect 1451 71 1453 75
rect 1457 71 1461 75
rect 1451 69 1461 71
rect 1464 75 1476 77
rect 1464 71 1468 75
rect 1472 71 1476 75
rect 1464 69 1476 71
rect 1479 75 1489 77
rect 1479 71 1483 75
rect 1487 71 1489 75
rect 1479 69 1489 71
rect 1493 75 1503 77
rect 1493 71 1495 75
rect 1499 71 1503 75
rect 1493 69 1503 71
rect 1505 75 1515 77
rect 1505 71 1509 75
rect 1513 71 1515 75
rect 1505 69 1515 71
rect 1621 75 1631 77
rect 1621 71 1623 75
rect 1627 71 1631 75
rect 1621 69 1631 71
rect 1634 75 1646 77
rect 1634 71 1638 75
rect 1642 71 1646 75
rect 1634 69 1646 71
rect 1649 75 1659 77
rect 1649 71 1653 75
rect 1657 71 1659 75
rect 1649 69 1659 71
rect 1663 75 1673 77
rect 1663 71 1665 75
rect 1669 71 1673 75
rect 1663 69 1673 71
rect 1675 75 1685 77
rect 1675 71 1679 75
rect 1683 71 1685 75
rect 1675 69 1685 71
rect 1975 75 1985 77
rect 1975 71 1977 75
rect 1981 71 1985 75
rect 1975 69 1985 71
rect 1988 75 2000 77
rect 1988 71 1992 75
rect 1996 71 2000 75
rect 1988 69 2000 71
rect 2003 75 2013 77
rect 2003 71 2007 75
rect 2011 71 2013 75
rect 2003 69 2013 71
rect 2017 75 2027 77
rect 2017 71 2019 75
rect 2023 71 2027 75
rect 2017 69 2027 71
rect 2029 75 2039 77
rect 2029 71 2033 75
rect 2037 71 2039 75
rect 2029 69 2039 71
rect 998 -61 1008 -59
rect 998 -65 1000 -61
rect 1004 -65 1008 -61
rect 998 -67 1008 -65
rect 1011 -61 1023 -59
rect 1011 -65 1015 -61
rect 1019 -65 1023 -61
rect 1011 -67 1023 -65
rect 1026 -61 1036 -59
rect 1026 -65 1030 -61
rect 1034 -65 1036 -61
rect 1026 -67 1036 -65
rect 931 -100 941 -98
rect 931 -104 933 -100
rect 937 -104 941 -100
rect 931 -106 941 -104
rect 944 -100 956 -98
rect 944 -104 948 -100
rect 952 -104 956 -100
rect 944 -106 956 -104
rect 959 -100 969 -98
rect 1066 -96 1076 -94
rect 959 -104 963 -100
rect 967 -104 969 -100
rect 959 -106 969 -104
rect 1066 -100 1068 -96
rect 1072 -100 1076 -96
rect 1066 -102 1076 -100
rect 1079 -96 1091 -94
rect 1079 -100 1083 -96
rect 1087 -100 1091 -96
rect 1079 -102 1091 -100
rect 1094 -96 1104 -94
rect 1094 -100 1098 -96
rect 1102 -100 1104 -96
rect 1094 -102 1104 -100
rect 998 -144 1008 -142
rect 998 -148 1000 -144
rect 1004 -148 1008 -144
rect 998 -150 1008 -148
rect 1011 -144 1023 -142
rect 1011 -148 1015 -144
rect 1019 -148 1023 -144
rect 1011 -150 1023 -148
rect 1026 -144 1036 -142
rect 1026 -148 1030 -144
rect 1034 -148 1036 -144
rect 1026 -150 1036 -148
rect 752 -245 762 -243
rect 752 -249 754 -245
rect 758 -249 762 -245
rect 752 -251 762 -249
rect 765 -245 777 -243
rect 765 -249 769 -245
rect 773 -249 777 -245
rect 765 -251 777 -249
rect 780 -245 790 -243
rect 780 -249 784 -245
rect 788 -249 790 -245
rect 780 -251 790 -249
rect 987 -245 997 -243
rect 987 -249 989 -245
rect 993 -249 997 -245
rect 987 -251 997 -249
rect 1000 -245 1012 -243
rect 1000 -249 1004 -245
rect 1008 -249 1012 -245
rect 1000 -251 1012 -249
rect 1015 -245 1025 -243
rect 1015 -249 1019 -245
rect 1023 -249 1025 -245
rect 1015 -251 1025 -249
rect 685 -284 695 -282
rect 685 -288 687 -284
rect 691 -288 695 -284
rect 685 -290 695 -288
rect 698 -284 710 -282
rect 698 -288 702 -284
rect 706 -288 710 -284
rect 698 -290 710 -288
rect 713 -284 723 -282
rect 820 -280 830 -278
rect 713 -288 717 -284
rect 721 -288 723 -284
rect 713 -290 723 -288
rect 820 -284 822 -280
rect 826 -284 830 -280
rect 820 -286 830 -284
rect 833 -280 845 -278
rect 833 -284 837 -280
rect 841 -284 845 -280
rect 833 -286 845 -284
rect 848 -280 858 -278
rect 848 -284 852 -280
rect 856 -284 858 -280
rect 848 -286 858 -284
rect 920 -284 930 -282
rect 920 -288 922 -284
rect 926 -288 930 -284
rect 920 -290 930 -288
rect 933 -284 945 -282
rect 933 -288 937 -284
rect 941 -288 945 -284
rect 933 -290 945 -288
rect 948 -284 958 -282
rect 1055 -280 1065 -278
rect 948 -288 952 -284
rect 956 -288 958 -284
rect 948 -290 958 -288
rect 752 -328 762 -326
rect 752 -332 754 -328
rect 758 -332 762 -328
rect 752 -334 762 -332
rect 765 -328 777 -326
rect 765 -332 769 -328
rect 773 -332 777 -328
rect 765 -334 777 -332
rect 780 -328 790 -326
rect 780 -332 784 -328
rect 788 -332 790 -328
rect 780 -334 790 -332
rect 666 -418 676 -416
rect 666 -422 668 -418
rect 672 -422 676 -418
rect 666 -424 676 -422
rect 679 -418 691 -416
rect 679 -422 683 -418
rect 687 -422 691 -418
rect 679 -424 691 -422
rect 694 -418 704 -416
rect 694 -422 698 -418
rect 702 -422 704 -418
rect 694 -424 704 -422
rect 708 -418 718 -416
rect 708 -422 710 -418
rect 714 -422 718 -418
rect 708 -424 718 -422
rect 720 -418 730 -416
rect 720 -422 724 -418
rect 728 -422 730 -418
rect 720 -424 730 -422
rect 1055 -284 1057 -280
rect 1061 -284 1065 -280
rect 1055 -286 1065 -284
rect 1068 -280 1080 -278
rect 1068 -284 1072 -280
rect 1076 -284 1080 -280
rect 1068 -286 1080 -284
rect 1083 -280 1093 -278
rect 1083 -284 1087 -280
rect 1091 -284 1093 -280
rect 1083 -286 1093 -284
rect 987 -328 997 -326
rect 987 -332 989 -328
rect 993 -332 997 -328
rect 987 -334 997 -332
rect 1000 -328 1012 -326
rect 1000 -332 1004 -328
rect 1008 -332 1012 -328
rect 1000 -334 1012 -332
rect 1015 -328 1025 -326
rect 1015 -332 1019 -328
rect 1023 -332 1025 -328
rect 1015 -334 1025 -332
rect 918 -418 928 -416
rect 918 -422 920 -418
rect 924 -422 928 -418
rect 918 -424 928 -422
rect 931 -418 943 -416
rect 931 -422 935 -418
rect 939 -422 943 -418
rect 931 -424 943 -422
rect 946 -418 956 -416
rect 946 -422 950 -418
rect 954 -422 956 -418
rect 946 -424 956 -422
rect 960 -418 970 -416
rect 960 -422 962 -418
rect 966 -422 970 -418
rect 960 -424 970 -422
rect 972 -418 982 -416
rect 972 -422 976 -418
rect 980 -422 982 -418
rect 972 -424 982 -422
rect 1035 -418 1045 -416
rect 1035 -422 1037 -418
rect 1041 -422 1045 -418
rect 1035 -424 1045 -422
rect 1048 -424 1060 -416
rect 1063 -418 1073 -416
rect 1063 -422 1067 -418
rect 1071 -422 1073 -418
rect 1063 -424 1073 -422
rect 1077 -418 1087 -416
rect 1077 -422 1079 -418
rect 1083 -422 1087 -418
rect 1077 -424 1087 -422
rect 1089 -418 1099 -416
rect 1089 -422 1093 -418
rect 1097 -422 1099 -418
rect 1089 -424 1099 -422
rect 2145 75 2155 77
rect 2145 71 2147 75
rect 2151 71 2155 75
rect 2145 69 2155 71
rect 2158 75 2170 77
rect 2158 71 2162 75
rect 2166 71 2170 75
rect 2158 69 2170 71
rect 2173 75 2183 77
rect 2173 71 2177 75
rect 2181 71 2183 75
rect 2173 69 2183 71
rect 2187 75 2197 77
rect 2187 71 2189 75
rect 2193 71 2197 75
rect 2187 69 2197 71
rect 2199 75 2209 77
rect 2199 71 2203 75
rect 2207 71 2209 75
rect 2199 69 2209 71
rect 1504 -61 1514 -59
rect 1504 -65 1506 -61
rect 1510 -65 1514 -61
rect 1504 -67 1514 -65
rect 1517 -61 1529 -59
rect 1517 -65 1521 -61
rect 1525 -65 1529 -61
rect 1517 -67 1529 -65
rect 1532 -61 1542 -59
rect 1532 -65 1536 -61
rect 1540 -65 1542 -61
rect 1532 -67 1542 -65
rect 1437 -100 1447 -98
rect 1437 -104 1439 -100
rect 1443 -104 1447 -100
rect 1437 -106 1447 -104
rect 1450 -100 1462 -98
rect 1450 -104 1454 -100
rect 1458 -104 1462 -100
rect 1450 -106 1462 -104
rect 1465 -100 1475 -98
rect 1572 -96 1582 -94
rect 1465 -104 1469 -100
rect 1473 -104 1475 -100
rect 1465 -106 1475 -104
rect 1572 -100 1574 -96
rect 1578 -100 1582 -96
rect 1572 -102 1582 -100
rect 1585 -96 1597 -94
rect 1585 -100 1589 -96
rect 1593 -100 1597 -96
rect 1585 -102 1597 -100
rect 1600 -96 1610 -94
rect 1600 -100 1604 -96
rect 1608 -100 1610 -96
rect 1600 -102 1610 -100
rect 1504 -144 1514 -142
rect 1504 -148 1506 -144
rect 1510 -148 1514 -144
rect 1504 -150 1514 -148
rect 1517 -144 1529 -142
rect 1517 -148 1521 -144
rect 1525 -148 1529 -144
rect 1517 -150 1529 -148
rect 1532 -144 1542 -142
rect 1532 -148 1536 -144
rect 1540 -148 1542 -144
rect 1532 -150 1542 -148
rect 1275 -245 1285 -243
rect 1275 -249 1277 -245
rect 1281 -249 1285 -245
rect 1275 -251 1285 -249
rect 1288 -245 1300 -243
rect 1288 -249 1292 -245
rect 1296 -249 1300 -245
rect 1288 -251 1300 -249
rect 1303 -245 1313 -243
rect 1303 -249 1307 -245
rect 1311 -249 1313 -245
rect 1303 -251 1313 -249
rect 1510 -245 1520 -243
rect 1510 -249 1512 -245
rect 1516 -249 1520 -245
rect 1510 -251 1520 -249
rect 1523 -245 1535 -243
rect 1523 -249 1527 -245
rect 1531 -249 1535 -245
rect 1523 -251 1535 -249
rect 1538 -245 1548 -243
rect 1538 -249 1542 -245
rect 1546 -249 1548 -245
rect 1538 -251 1548 -249
rect 1208 -284 1218 -282
rect 1208 -288 1210 -284
rect 1214 -288 1218 -284
rect 1208 -290 1218 -288
rect 1221 -284 1233 -282
rect 1221 -288 1225 -284
rect 1229 -288 1233 -284
rect 1221 -290 1233 -288
rect 1236 -284 1246 -282
rect 1343 -280 1353 -278
rect 1236 -288 1240 -284
rect 1244 -288 1246 -284
rect 1236 -290 1246 -288
rect 1343 -284 1345 -280
rect 1349 -284 1353 -280
rect 1343 -286 1353 -284
rect 1356 -280 1368 -278
rect 1356 -284 1360 -280
rect 1364 -284 1368 -280
rect 1356 -286 1368 -284
rect 1371 -280 1381 -278
rect 1371 -284 1375 -280
rect 1379 -284 1381 -280
rect 1371 -286 1381 -284
rect 1443 -284 1453 -282
rect 1443 -288 1445 -284
rect 1449 -288 1453 -284
rect 1443 -290 1453 -288
rect 1456 -284 1468 -282
rect 1456 -288 1460 -284
rect 1464 -288 1468 -284
rect 1456 -290 1468 -288
rect 1471 -284 1481 -282
rect 1578 -280 1588 -278
rect 1471 -288 1475 -284
rect 1479 -288 1481 -284
rect 1471 -290 1481 -288
rect 1275 -328 1285 -326
rect 1275 -332 1277 -328
rect 1281 -332 1285 -328
rect 1275 -334 1285 -332
rect 1288 -328 1300 -326
rect 1288 -332 1292 -328
rect 1296 -332 1300 -328
rect 1288 -334 1300 -332
rect 1303 -328 1313 -326
rect 1303 -332 1307 -328
rect 1311 -332 1313 -328
rect 1303 -334 1313 -332
rect 1189 -418 1199 -416
rect 1189 -422 1191 -418
rect 1195 -422 1199 -418
rect 1189 -424 1199 -422
rect 1202 -418 1214 -416
rect 1202 -422 1206 -418
rect 1210 -422 1214 -418
rect 1202 -424 1214 -422
rect 1217 -418 1227 -416
rect 1217 -422 1221 -418
rect 1225 -422 1227 -418
rect 1217 -424 1227 -422
rect 1231 -418 1241 -416
rect 1231 -422 1233 -418
rect 1237 -422 1241 -418
rect 1231 -424 1241 -422
rect 1243 -418 1253 -416
rect 1243 -422 1247 -418
rect 1251 -422 1253 -418
rect 1243 -424 1253 -422
rect 1578 -284 1580 -280
rect 1584 -284 1588 -280
rect 1578 -286 1588 -284
rect 1591 -280 1603 -278
rect 1591 -284 1595 -280
rect 1599 -284 1603 -280
rect 1591 -286 1603 -284
rect 1606 -280 1616 -278
rect 1606 -284 1610 -280
rect 1614 -284 1616 -280
rect 1606 -286 1616 -284
rect 1510 -328 1520 -326
rect 1510 -332 1512 -328
rect 1516 -332 1520 -328
rect 1510 -334 1520 -332
rect 1523 -328 1535 -326
rect 1523 -332 1527 -328
rect 1531 -332 1535 -328
rect 1523 -334 1535 -332
rect 1538 -328 1548 -326
rect 1538 -332 1542 -328
rect 1546 -332 1548 -328
rect 1538 -334 1548 -332
rect 1441 -418 1451 -416
rect 1441 -422 1443 -418
rect 1447 -422 1451 -418
rect 1441 -424 1451 -422
rect 1454 -418 1466 -416
rect 1454 -422 1458 -418
rect 1462 -422 1466 -418
rect 1454 -424 1466 -422
rect 1469 -418 1479 -416
rect 1469 -422 1473 -418
rect 1477 -422 1479 -418
rect 1469 -424 1479 -422
rect 1483 -418 1493 -416
rect 1483 -422 1485 -418
rect 1489 -422 1493 -418
rect 1483 -424 1493 -422
rect 1495 -418 1505 -416
rect 1495 -422 1499 -418
rect 1503 -422 1505 -418
rect 1495 -424 1505 -422
rect 1558 -418 1568 -416
rect 1558 -422 1560 -418
rect 1564 -422 1568 -418
rect 1558 -424 1568 -422
rect 1571 -424 1583 -416
rect 1586 -418 1596 -416
rect 1586 -422 1590 -418
rect 1594 -422 1596 -418
rect 1586 -424 1596 -422
rect 1600 -418 1610 -416
rect 1600 -422 1602 -418
rect 1606 -422 1610 -418
rect 1600 -424 1610 -422
rect 1612 -418 1622 -416
rect 1612 -422 1616 -418
rect 1620 -422 1622 -418
rect 1612 -424 1622 -422
rect 2028 -61 2038 -59
rect 2028 -65 2030 -61
rect 2034 -65 2038 -61
rect 2028 -67 2038 -65
rect 2041 -61 2053 -59
rect 2041 -65 2045 -61
rect 2049 -65 2053 -61
rect 2041 -67 2053 -65
rect 2056 -61 2066 -59
rect 2056 -65 2060 -61
rect 2064 -65 2066 -61
rect 2056 -67 2066 -65
rect 1961 -100 1971 -98
rect 1961 -104 1963 -100
rect 1967 -104 1971 -100
rect 1961 -106 1971 -104
rect 1974 -100 1986 -98
rect 1974 -104 1978 -100
rect 1982 -104 1986 -100
rect 1974 -106 1986 -104
rect 1989 -100 1999 -98
rect 2096 -96 2106 -94
rect 1989 -104 1993 -100
rect 1997 -104 1999 -100
rect 1989 -106 1999 -104
rect 2096 -100 2098 -96
rect 2102 -100 2106 -96
rect 2096 -102 2106 -100
rect 2109 -96 2121 -94
rect 2109 -100 2113 -96
rect 2117 -100 2121 -96
rect 2109 -102 2121 -100
rect 2124 -96 2134 -94
rect 2124 -100 2128 -96
rect 2132 -100 2134 -96
rect 2124 -102 2134 -100
rect 2028 -144 2038 -142
rect 2028 -148 2030 -144
rect 2034 -148 2038 -144
rect 2028 -150 2038 -148
rect 2041 -144 2053 -142
rect 2041 -148 2045 -144
rect 2049 -148 2053 -144
rect 2041 -150 2053 -148
rect 2056 -144 2066 -142
rect 2056 -148 2060 -144
rect 2064 -148 2066 -144
rect 2056 -150 2066 -148
rect 1798 -245 1808 -243
rect 1798 -249 1800 -245
rect 1804 -249 1808 -245
rect 1798 -251 1808 -249
rect 1811 -245 1823 -243
rect 1811 -249 1815 -245
rect 1819 -249 1823 -245
rect 1811 -251 1823 -249
rect 1826 -245 1836 -243
rect 1826 -249 1830 -245
rect 1834 -249 1836 -245
rect 1826 -251 1836 -249
rect 2033 -245 2043 -243
rect 2033 -249 2035 -245
rect 2039 -249 2043 -245
rect 2033 -251 2043 -249
rect 2046 -245 2058 -243
rect 2046 -249 2050 -245
rect 2054 -249 2058 -245
rect 2046 -251 2058 -249
rect 2061 -245 2071 -243
rect 2061 -249 2065 -245
rect 2069 -249 2071 -245
rect 2061 -251 2071 -249
rect 1731 -284 1741 -282
rect 1731 -288 1733 -284
rect 1737 -288 1741 -284
rect 1731 -290 1741 -288
rect 1744 -284 1756 -282
rect 1744 -288 1748 -284
rect 1752 -288 1756 -284
rect 1744 -290 1756 -288
rect 1759 -284 1769 -282
rect 1866 -280 1876 -278
rect 1759 -288 1763 -284
rect 1767 -288 1769 -284
rect 1759 -290 1769 -288
rect 1866 -284 1868 -280
rect 1872 -284 1876 -280
rect 1866 -286 1876 -284
rect 1879 -280 1891 -278
rect 1879 -284 1883 -280
rect 1887 -284 1891 -280
rect 1879 -286 1891 -284
rect 1894 -280 1904 -278
rect 1894 -284 1898 -280
rect 1902 -284 1904 -280
rect 1894 -286 1904 -284
rect 1966 -284 1976 -282
rect 1966 -288 1968 -284
rect 1972 -288 1976 -284
rect 1966 -290 1976 -288
rect 1979 -284 1991 -282
rect 1979 -288 1983 -284
rect 1987 -288 1991 -284
rect 1979 -290 1991 -288
rect 1994 -284 2004 -282
rect 2101 -280 2111 -278
rect 1994 -288 1998 -284
rect 2002 -288 2004 -284
rect 1994 -290 2004 -288
rect 1798 -328 1808 -326
rect 1798 -332 1800 -328
rect 1804 -332 1808 -328
rect 1798 -334 1808 -332
rect 1811 -328 1823 -326
rect 1811 -332 1815 -328
rect 1819 -332 1823 -328
rect 1811 -334 1823 -332
rect 1826 -328 1836 -326
rect 1826 -332 1830 -328
rect 1834 -332 1836 -328
rect 1826 -334 1836 -332
rect 1712 -418 1722 -416
rect 1712 -422 1714 -418
rect 1718 -422 1722 -418
rect 1712 -424 1722 -422
rect 1725 -418 1737 -416
rect 1725 -422 1729 -418
rect 1733 -422 1737 -418
rect 1725 -424 1737 -422
rect 1740 -418 1750 -416
rect 1740 -422 1744 -418
rect 1748 -422 1750 -418
rect 1740 -424 1750 -422
rect 1754 -418 1764 -416
rect 1754 -422 1756 -418
rect 1760 -422 1764 -418
rect 1754 -424 1764 -422
rect 1766 -418 1776 -416
rect 1766 -422 1770 -418
rect 1774 -422 1776 -418
rect 1766 -424 1776 -422
rect 2101 -284 2103 -280
rect 2107 -284 2111 -280
rect 2101 -286 2111 -284
rect 2114 -280 2126 -278
rect 2114 -284 2118 -280
rect 2122 -284 2126 -280
rect 2114 -286 2126 -284
rect 2129 -280 2139 -278
rect 2129 -284 2133 -280
rect 2137 -284 2139 -280
rect 2129 -286 2139 -284
rect 2033 -328 2043 -326
rect 2033 -332 2035 -328
rect 2039 -332 2043 -328
rect 2033 -334 2043 -332
rect 2046 -328 2058 -326
rect 2046 -332 2050 -328
rect 2054 -332 2058 -328
rect 2046 -334 2058 -332
rect 2061 -328 2071 -326
rect 2061 -332 2065 -328
rect 2069 -332 2071 -328
rect 2061 -334 2071 -332
rect 1964 -418 1974 -416
rect 1964 -422 1966 -418
rect 1970 -422 1974 -418
rect 1964 -424 1974 -422
rect 1977 -418 1989 -416
rect 1977 -422 1981 -418
rect 1985 -422 1989 -418
rect 1977 -424 1989 -422
rect 1992 -418 2002 -416
rect 1992 -422 1996 -418
rect 2000 -422 2002 -418
rect 1992 -424 2002 -422
rect 2006 -418 2016 -416
rect 2006 -422 2008 -418
rect 2012 -422 2016 -418
rect 2006 -424 2016 -422
rect 2018 -418 2028 -416
rect 2018 -422 2022 -418
rect 2026 -422 2028 -418
rect 2018 -424 2028 -422
rect 2081 -418 2091 -416
rect 2081 -422 2083 -418
rect 2087 -422 2091 -418
rect 2081 -424 2091 -422
rect 2094 -424 2106 -416
rect 2109 -418 2119 -416
rect 2109 -422 2113 -418
rect 2117 -422 2119 -418
rect 2109 -424 2119 -422
rect 2123 -418 2133 -416
rect 2123 -422 2125 -418
rect 2129 -422 2133 -418
rect 2123 -424 2133 -422
rect 2135 -418 2145 -416
rect 2135 -422 2139 -418
rect 2143 -422 2145 -418
rect 2135 -424 2145 -422
rect 2321 -245 2331 -243
rect 2321 -249 2323 -245
rect 2327 -249 2331 -245
rect 2321 -251 2331 -249
rect 2334 -245 2346 -243
rect 2334 -249 2338 -245
rect 2342 -249 2346 -245
rect 2334 -251 2346 -249
rect 2349 -245 2359 -243
rect 2349 -249 2353 -245
rect 2357 -249 2359 -245
rect 2349 -251 2359 -249
rect 2556 -245 2566 -243
rect 2556 -249 2558 -245
rect 2562 -249 2566 -245
rect 2556 -251 2566 -249
rect 2569 -245 2581 -243
rect 2569 -249 2573 -245
rect 2577 -249 2581 -245
rect 2569 -251 2581 -249
rect 2584 -245 2594 -243
rect 2584 -249 2588 -245
rect 2592 -249 2594 -245
rect 2584 -251 2594 -249
rect 2254 -284 2264 -282
rect 2254 -288 2256 -284
rect 2260 -288 2264 -284
rect 2254 -290 2264 -288
rect 2267 -284 2279 -282
rect 2267 -288 2271 -284
rect 2275 -288 2279 -284
rect 2267 -290 2279 -288
rect 2282 -284 2292 -282
rect 2389 -280 2399 -278
rect 2282 -288 2286 -284
rect 2290 -288 2292 -284
rect 2282 -290 2292 -288
rect 2389 -284 2391 -280
rect 2395 -284 2399 -280
rect 2389 -286 2399 -284
rect 2402 -280 2414 -278
rect 2402 -284 2406 -280
rect 2410 -284 2414 -280
rect 2402 -286 2414 -284
rect 2417 -280 2427 -278
rect 2417 -284 2421 -280
rect 2425 -284 2427 -280
rect 2417 -286 2427 -284
rect 2489 -284 2499 -282
rect 2489 -288 2491 -284
rect 2495 -288 2499 -284
rect 2489 -290 2499 -288
rect 2502 -284 2514 -282
rect 2502 -288 2506 -284
rect 2510 -288 2514 -284
rect 2502 -290 2514 -288
rect 2517 -284 2527 -282
rect 2624 -280 2634 -278
rect 2517 -288 2521 -284
rect 2525 -288 2527 -284
rect 2517 -290 2527 -288
rect 2321 -328 2331 -326
rect 2321 -332 2323 -328
rect 2327 -332 2331 -328
rect 2321 -334 2331 -332
rect 2334 -328 2346 -326
rect 2334 -332 2338 -328
rect 2342 -332 2346 -328
rect 2334 -334 2346 -332
rect 2349 -328 2359 -326
rect 2349 -332 2353 -328
rect 2357 -332 2359 -328
rect 2349 -334 2359 -332
rect 2235 -418 2245 -416
rect 2235 -422 2237 -418
rect 2241 -422 2245 -418
rect 2235 -424 2245 -422
rect 2248 -418 2260 -416
rect 2248 -422 2252 -418
rect 2256 -422 2260 -418
rect 2248 -424 2260 -422
rect 2263 -418 2273 -416
rect 2263 -422 2267 -418
rect 2271 -422 2273 -418
rect 2263 -424 2273 -422
rect 2277 -418 2287 -416
rect 2277 -422 2279 -418
rect 2283 -422 2287 -418
rect 2277 -424 2287 -422
rect 2289 -418 2299 -416
rect 2289 -422 2293 -418
rect 2297 -422 2299 -418
rect 2289 -424 2299 -422
rect 2624 -284 2626 -280
rect 2630 -284 2634 -280
rect 2624 -286 2634 -284
rect 2637 -280 2649 -278
rect 2637 -284 2641 -280
rect 2645 -284 2649 -280
rect 2637 -286 2649 -284
rect 2652 -280 2662 -278
rect 2652 -284 2656 -280
rect 2660 -284 2662 -280
rect 2652 -286 2662 -284
rect 2556 -328 2566 -326
rect 2556 -332 2558 -328
rect 2562 -332 2566 -328
rect 2556 -334 2566 -332
rect 2569 -328 2581 -326
rect 2569 -332 2573 -328
rect 2577 -332 2581 -328
rect 2569 -334 2581 -332
rect 2584 -328 2594 -326
rect 2584 -332 2588 -328
rect 2592 -332 2594 -328
rect 2584 -334 2594 -332
rect 2487 -418 2497 -416
rect 2487 -422 2489 -418
rect 2493 -422 2497 -418
rect 2487 -424 2497 -422
rect 2500 -418 2512 -416
rect 2500 -422 2504 -418
rect 2508 -422 2512 -418
rect 2500 -424 2512 -422
rect 2515 -418 2525 -416
rect 2515 -422 2519 -418
rect 2523 -422 2525 -418
rect 2515 -424 2525 -422
rect 2529 -418 2539 -416
rect 2529 -422 2531 -418
rect 2535 -422 2539 -418
rect 2529 -424 2539 -422
rect 2541 -418 2551 -416
rect 2541 -422 2545 -418
rect 2549 -422 2551 -418
rect 2541 -424 2551 -422
rect 2604 -418 2614 -416
rect 2604 -422 2606 -418
rect 2610 -422 2614 -418
rect 2604 -424 2614 -422
rect 2617 -424 2629 -416
rect 2632 -418 2642 -416
rect 2632 -422 2636 -418
rect 2640 -422 2642 -418
rect 2632 -424 2642 -422
rect 2646 -418 2656 -416
rect 2646 -422 2648 -418
rect 2652 -422 2656 -418
rect 2646 -424 2656 -422
rect 2658 -418 2668 -416
rect 2658 -422 2662 -418
rect 2666 -422 2668 -418
rect 2658 -424 2668 -422
<< metal1 >>
rect 81 1540 85 1576
rect 6 1536 9 1540
rect 13 1536 24 1540
rect 28 1536 40 1540
rect 44 1536 70 1540
rect 74 1536 96 1540
rect 100 1536 120 1540
rect 124 1536 131 1540
rect 24 1528 28 1536
rect 51 1528 55 1536
rect 75 1528 79 1536
rect 101 1528 105 1536
rect 125 1528 129 1536
rect 10 1506 14 1524
rect 36 1508 40 1524
rect 61 1519 65 1524
rect 87 1519 91 1524
rect 111 1519 115 1524
rect 61 1515 115 1519
rect 125 1515 1290 1519
rect 61 1508 65 1515
rect 101 1508 880 1512
rect 6 1502 14 1506
rect 24 1504 65 1508
rect 10 1487 14 1502
rect 36 1487 40 1504
rect 75 1501 526 1505
rect 51 1494 173 1498
rect 24 1473 28 1483
rect 125 1473 129 1483
rect 6 1469 10 1473
rect 14 1469 24 1473
rect 28 1469 42 1473
rect 46 1469 70 1473
rect 74 1469 96 1473
rect 100 1469 120 1473
rect 124 1469 133 1473
rect 55 1272 59 1469
rect 168 1306 173 1494
rect 231 1372 235 1398
rect 246 1372 250 1389
rect 489 1381 491 1385
rect 196 1335 197 1339
rect 201 1335 212 1339
rect 216 1335 228 1339
rect 232 1335 279 1339
rect 283 1338 295 1339
rect 283 1335 304 1338
rect 212 1327 216 1335
rect 284 1327 288 1335
rect 292 1334 304 1335
rect 308 1334 319 1338
rect 323 1334 335 1338
rect 339 1334 356 1338
rect 360 1334 372 1338
rect 376 1334 387 1338
rect 391 1334 393 1338
rect 319 1326 323 1334
rect 361 1326 365 1334
rect 387 1326 391 1334
rect 198 1306 202 1323
rect 224 1308 228 1323
rect 168 1302 202 1306
rect 212 1304 228 1308
rect 305 1305 309 1322
rect 331 1307 335 1322
rect 373 1315 377 1322
rect 362 1311 377 1315
rect 387 1312 393 1316
rect 198 1286 202 1302
rect 224 1297 228 1304
rect 297 1301 309 1305
rect 319 1303 335 1307
rect 347 1303 362 1307
rect 297 1297 301 1301
rect 224 1293 273 1297
rect 284 1293 301 1297
rect 239 1286 243 1293
rect 212 1272 216 1282
rect 254 1286 258 1293
rect 269 1286 273 1293
rect 305 1286 309 1301
rect 331 1299 335 1303
rect 358 1299 362 1303
rect 331 1295 350 1299
rect 358 1295 363 1299
rect 346 1286 350 1295
rect 373 1286 377 1311
rect 431 1299 435 1338
rect 448 1316 452 1338
rect 450 1312 452 1316
rect 388 1295 393 1299
rect 433 1295 435 1299
rect 224 1272 228 1282
rect 284 1272 288 1282
rect 319 1272 323 1282
rect 331 1272 335 1282
rect 361 1272 365 1282
rect 387 1272 391 1282
rect 55 1268 198 1272
rect 202 1268 212 1272
rect 216 1268 230 1272
rect 234 1268 279 1272
rect 283 1268 305 1272
rect 309 1268 319 1272
rect 323 1268 337 1272
rect 341 1268 356 1272
rect 360 1268 373 1272
rect 377 1268 387 1272
rect 391 1268 395 1272
rect 55 1067 59 1268
rect 303 1193 307 1197
rect 288 1189 292 1193
rect 296 1189 313 1193
rect 317 1189 322 1193
rect 318 1181 322 1189
rect 288 1162 292 1177
rect 319 1166 349 1170
rect 272 1158 292 1162
rect 304 1158 339 1162
rect 183 1149 224 1153
rect 183 1136 187 1149
rect 220 1141 224 1149
rect 228 1141 245 1145
rect 249 1141 254 1145
rect 159 1132 162 1136
rect 166 1132 177 1136
rect 181 1132 187 1136
rect 250 1133 254 1141
rect 177 1124 181 1132
rect 163 1113 167 1120
rect 220 1114 224 1129
rect 272 1122 276 1158
rect 288 1154 292 1158
rect 288 1150 307 1154
rect 303 1141 307 1150
rect 288 1127 292 1137
rect 318 1127 322 1137
rect 286 1123 294 1127
rect 298 1123 313 1127
rect 317 1123 323 1127
rect 251 1118 276 1122
rect 335 1118 339 1158
rect 344 1157 349 1166
rect 344 1153 399 1157
rect 354 1145 359 1149
rect 363 1145 380 1149
rect 384 1145 391 1149
rect 385 1137 389 1145
rect 355 1118 359 1133
rect 394 1126 399 1153
rect 431 1126 435 1295
rect 386 1122 410 1126
rect 433 1122 435 1126
rect 335 1114 359 1118
rect 371 1114 410 1118
rect 157 1109 167 1113
rect 177 1110 224 1114
rect 236 1110 276 1114
rect 163 1102 167 1109
rect 220 1106 224 1110
rect 220 1102 239 1106
rect 177 1088 181 1098
rect 235 1093 239 1102
rect 159 1084 163 1088
rect 167 1084 177 1088
rect 181 1084 189 1088
rect 185 1079 189 1084
rect 220 1079 224 1089
rect 250 1079 254 1089
rect 272 1079 276 1110
rect 288 1106 292 1110
rect 296 1106 313 1110
rect 317 1106 324 1110
rect 318 1098 322 1106
rect 288 1079 292 1094
rect 335 1087 339 1114
rect 355 1110 359 1114
rect 355 1106 374 1110
rect 370 1097 374 1106
rect 319 1083 339 1087
rect 355 1083 359 1093
rect 385 1083 389 1093
rect 356 1079 361 1083
rect 365 1079 380 1083
rect 384 1079 393 1083
rect 185 1075 226 1079
rect 230 1075 245 1079
rect 249 1075 256 1079
rect 272 1075 292 1079
rect 304 1075 330 1079
rect 396 1075 401 1114
rect 288 1071 292 1075
rect 326 1071 401 1075
rect 288 1067 307 1071
rect 55 1063 156 1067
rect -97 1037 -96 1041
rect -92 1037 -81 1041
rect -77 1037 -65 1041
rect -61 1037 -14 1041
rect -10 1037 -3 1041
rect -81 1029 -77 1037
rect -9 1029 -5 1037
rect -95 1008 -91 1025
rect -69 1010 -65 1025
rect -54 1016 -1 1020
rect -99 1004 -91 1008
rect -81 1006 -65 1010
rect -39 1009 -1 1013
rect -95 988 -91 1004
rect -69 999 -65 1006
rect -24 1002 -1 1006
rect -69 995 -20 999
rect -9 995 -1 999
rect -54 988 -50 995
rect -81 974 -77 984
rect -39 988 -35 995
rect -24 988 -20 995
rect -69 974 -65 984
rect -9 974 -5 984
rect -99 970 -95 974
rect -91 970 -81 974
rect -77 970 -63 974
rect -59 970 -14 974
rect -10 970 -3 974
rect -42 959 -38 970
rect 55 959 59 1063
rect 152 1044 156 1063
rect 303 1058 307 1067
rect 288 1044 292 1054
rect 318 1044 322 1054
rect 152 1040 294 1044
rect 298 1040 313 1044
rect 317 1040 324 1044
rect 222 985 226 1008
rect 232 985 236 999
rect 182 964 183 968
rect 187 964 198 968
rect 202 964 214 968
rect 218 964 265 968
rect 269 967 281 968
rect 269 964 290 967
rect -42 955 59 959
rect 198 956 202 964
rect 270 956 274 964
rect 278 963 290 964
rect 294 963 305 967
rect 309 963 321 967
rect 325 963 342 967
rect 346 963 358 967
rect 362 963 373 967
rect 377 963 379 967
rect 305 955 309 963
rect 347 955 351 963
rect 373 955 377 963
rect 184 935 188 952
rect 210 937 214 952
rect 140 931 188 935
rect 198 933 214 937
rect 291 934 295 951
rect 317 936 321 951
rect 359 944 363 951
rect 431 945 435 1122
rect 448 1118 452 1312
rect 450 1114 452 1118
rect 348 940 363 944
rect 373 941 379 945
rect 433 941 435 945
rect -45 873 -44 877
rect -40 873 -29 877
rect -25 873 -13 877
rect -9 873 17 877
rect 21 873 43 877
rect 47 873 67 877
rect 71 873 78 877
rect -29 865 -25 873
rect -2 865 2 873
rect 22 865 26 873
rect 48 865 52 873
rect 72 865 76 873
rect -43 843 -39 861
rect -17 845 -13 861
rect 8 856 12 861
rect 34 856 38 861
rect 58 856 62 861
rect 140 856 144 931
rect 184 915 188 931
rect 210 926 214 933
rect 283 930 295 934
rect 305 932 321 936
rect 333 932 348 936
rect 283 926 287 930
rect 210 922 259 926
rect 270 922 287 926
rect 225 915 229 922
rect 198 901 202 911
rect 240 915 244 922
rect 255 915 259 922
rect 291 915 295 930
rect 317 928 321 932
rect 344 928 348 932
rect 317 924 336 928
rect 344 924 349 928
rect 332 915 336 924
rect 359 915 363 940
rect 374 924 379 928
rect 210 901 214 911
rect 270 901 274 911
rect 305 901 309 911
rect 317 901 321 911
rect 347 901 351 911
rect 373 901 377 911
rect 182 897 184 901
rect 188 897 198 901
rect 202 897 216 901
rect 220 897 265 901
rect 269 897 291 901
rect 295 897 305 901
rect 309 897 323 901
rect 327 897 342 901
rect 346 897 359 901
rect 363 897 373 901
rect 377 897 379 901
rect 8 852 62 856
rect 72 852 144 856
rect 8 845 12 852
rect 431 849 435 941
rect 448 928 452 1114
rect 487 1121 491 1381
rect 522 1308 526 1501
rect 588 1382 592 1398
rect 835 1391 838 1395
rect 552 1337 554 1341
rect 558 1337 569 1341
rect 573 1337 585 1341
rect 589 1337 621 1341
rect 625 1340 641 1341
rect 625 1337 650 1340
rect 569 1329 573 1337
rect 626 1329 630 1337
rect 636 1336 650 1337
rect 654 1336 665 1340
rect 669 1336 681 1340
rect 685 1336 702 1340
rect 706 1336 718 1340
rect 722 1336 733 1340
rect 737 1336 739 1340
rect 665 1328 669 1336
rect 707 1328 711 1336
rect 733 1328 737 1336
rect 555 1308 559 1325
rect 581 1310 585 1325
rect 596 1316 636 1320
rect 522 1304 559 1308
rect 569 1306 585 1310
rect 651 1307 655 1324
rect 677 1309 681 1324
rect 719 1317 723 1324
rect 708 1313 723 1317
rect 733 1314 739 1318
rect 555 1288 559 1304
rect 581 1299 585 1306
rect 641 1303 655 1307
rect 665 1305 681 1309
rect 693 1305 708 1309
rect 641 1299 645 1303
rect 581 1295 615 1299
rect 626 1295 645 1299
rect 596 1288 600 1295
rect 569 1274 573 1284
rect 611 1288 615 1295
rect 651 1288 655 1303
rect 677 1301 681 1305
rect 704 1301 708 1305
rect 677 1297 696 1301
rect 704 1297 709 1301
rect 692 1288 696 1297
rect 719 1288 723 1313
rect 775 1301 779 1361
rect 792 1318 796 1370
rect 794 1314 796 1318
rect 734 1297 739 1301
rect 777 1297 779 1301
rect 581 1274 585 1284
rect 626 1274 630 1284
rect 665 1274 669 1284
rect 677 1274 681 1284
rect 707 1274 711 1284
rect 733 1274 737 1284
rect 551 1270 555 1274
rect 559 1270 569 1274
rect 573 1270 587 1274
rect 591 1270 621 1274
rect 625 1270 651 1274
rect 655 1270 665 1274
rect 669 1270 683 1274
rect 687 1270 702 1274
rect 706 1270 719 1274
rect 723 1270 733 1274
rect 737 1270 740 1274
rect 647 1201 651 1205
rect 632 1197 636 1201
rect 640 1197 657 1201
rect 661 1197 666 1201
rect 662 1189 666 1197
rect 632 1170 636 1185
rect 663 1174 693 1178
rect 616 1166 636 1170
rect 648 1166 683 1170
rect 527 1157 568 1161
rect 527 1144 531 1157
rect 564 1149 568 1157
rect 572 1149 589 1153
rect 593 1149 598 1153
rect 503 1140 506 1144
rect 510 1140 521 1144
rect 525 1140 531 1144
rect 594 1141 598 1149
rect 521 1132 525 1140
rect 507 1121 511 1128
rect 564 1122 568 1137
rect 616 1130 620 1166
rect 632 1162 636 1166
rect 632 1158 651 1162
rect 647 1149 651 1158
rect 632 1135 636 1145
rect 662 1135 666 1145
rect 630 1131 638 1135
rect 642 1131 657 1135
rect 661 1131 667 1135
rect 595 1126 620 1130
rect 679 1126 683 1166
rect 688 1165 693 1174
rect 688 1161 743 1165
rect 698 1153 703 1157
rect 707 1153 724 1157
rect 728 1153 735 1157
rect 729 1145 733 1153
rect 699 1126 703 1141
rect 738 1134 743 1161
rect 775 1134 779 1297
rect 730 1130 754 1134
rect 777 1130 779 1134
rect 679 1122 703 1126
rect 715 1122 754 1126
rect 487 1117 511 1121
rect 521 1118 568 1122
rect 580 1118 620 1122
rect 487 1014 491 1117
rect 507 1110 511 1117
rect 564 1114 568 1118
rect 564 1110 583 1114
rect 521 1096 525 1106
rect 579 1101 583 1110
rect 503 1092 507 1096
rect 511 1092 521 1096
rect 525 1092 533 1096
rect 529 1087 533 1092
rect 564 1087 568 1097
rect 594 1087 598 1097
rect 616 1087 620 1118
rect 632 1114 636 1118
rect 640 1114 657 1118
rect 661 1114 668 1118
rect 662 1106 666 1114
rect 632 1087 636 1102
rect 679 1095 683 1122
rect 699 1118 703 1122
rect 699 1114 718 1118
rect 714 1105 718 1114
rect 663 1091 683 1095
rect 699 1091 703 1101
rect 729 1091 733 1101
rect 700 1087 705 1091
rect 709 1087 724 1091
rect 728 1087 737 1091
rect 529 1083 570 1087
rect 574 1083 589 1087
rect 593 1083 600 1087
rect 616 1083 636 1087
rect 648 1083 674 1087
rect 740 1083 745 1122
rect 632 1079 636 1083
rect 670 1079 745 1083
rect 632 1075 651 1079
rect 647 1066 651 1075
rect 632 1052 636 1062
rect 662 1052 666 1062
rect 630 1048 638 1052
rect 642 1048 657 1052
rect 661 1048 668 1052
rect 489 1010 491 1014
rect 564 983 568 999
rect 525 972 526 976
rect 530 972 541 976
rect 545 972 557 976
rect 561 972 593 976
rect 597 975 613 976
rect 597 972 622 975
rect 541 964 545 972
rect 598 964 602 972
rect 608 971 622 972
rect 626 971 637 975
rect 641 971 653 975
rect 657 971 674 975
rect 678 971 690 975
rect 694 971 705 975
rect 709 971 711 975
rect 637 963 641 971
rect 679 963 683 971
rect 705 963 709 971
rect 527 943 531 960
rect 553 945 557 960
rect 568 951 608 955
rect 450 924 452 928
rect 448 849 452 924
rect 506 939 531 943
rect 541 941 557 945
rect 623 942 627 959
rect 649 944 653 959
rect 691 952 695 959
rect 775 953 779 1130
rect 792 1126 796 1314
rect 794 1122 796 1126
rect 680 948 695 952
rect 705 949 711 953
rect 777 949 779 953
rect 506 849 510 939
rect 527 923 531 939
rect 553 934 557 941
rect 613 938 627 942
rect 637 940 653 944
rect 665 940 680 944
rect 613 934 617 938
rect 553 930 587 934
rect 598 930 617 934
rect 568 923 572 930
rect 541 909 545 919
rect 583 923 587 930
rect 623 923 627 938
rect 649 936 653 940
rect 676 936 680 940
rect 649 932 668 936
rect 676 932 681 936
rect 664 923 668 932
rect 691 923 695 948
rect 706 932 711 936
rect 553 909 557 919
rect 598 909 602 919
rect 637 909 641 919
rect 649 909 653 919
rect 679 909 683 919
rect 705 909 709 919
rect 525 905 527 909
rect 531 905 541 909
rect 545 905 559 909
rect 563 905 593 909
rect 597 905 623 909
rect 627 905 637 909
rect 641 905 655 909
rect 659 905 674 909
rect 678 905 691 909
rect 695 905 705 909
rect 709 905 712 909
rect 48 845 133 849
rect 508 845 510 849
rect -47 839 -39 843
rect -29 841 12 845
rect 431 842 435 845
rect 448 842 452 845
rect 775 842 779 949
rect 792 936 796 1122
rect 833 1126 838 1391
rect 876 1322 880 1508
rect 1178 1400 1184 1404
rect 895 1351 898 1355
rect 902 1351 913 1355
rect 917 1351 929 1355
rect 933 1351 950 1355
rect 954 1351 975 1355
rect 979 1351 990 1355
rect 994 1351 1006 1355
rect 1010 1351 1027 1355
rect 1031 1351 1043 1355
rect 1047 1351 1058 1355
rect 1062 1351 1064 1355
rect 913 1343 917 1351
rect 955 1343 959 1351
rect 990 1343 994 1351
rect 1032 1343 1036 1351
rect 1058 1343 1062 1351
rect 899 1322 903 1339
rect 925 1324 929 1339
rect 976 1324 980 1339
rect 1002 1324 1006 1339
rect 1044 1332 1048 1339
rect 1033 1328 1048 1332
rect 1058 1329 1064 1333
rect 876 1318 903 1322
rect 913 1320 929 1324
rect 941 1320 980 1324
rect 990 1320 1006 1324
rect 1018 1320 1033 1324
rect 899 1303 903 1318
rect 925 1316 929 1320
rect 925 1312 944 1316
rect 940 1303 944 1312
rect 976 1303 980 1320
rect 1002 1316 1006 1320
rect 1029 1316 1033 1320
rect 1002 1312 1021 1316
rect 1029 1312 1034 1316
rect 1017 1303 1021 1312
rect 1044 1303 1048 1328
rect 1133 1316 1137 1355
rect 1150 1333 1154 1355
rect 1152 1329 1154 1333
rect 1059 1312 1064 1316
rect 1135 1312 1137 1316
rect 913 1289 917 1299
rect 925 1289 929 1299
rect 955 1289 959 1299
rect 990 1289 994 1299
rect 1002 1289 1006 1299
rect 1032 1289 1036 1299
rect 1058 1289 1062 1299
rect 898 1285 899 1289
rect 903 1285 913 1289
rect 917 1285 931 1289
rect 935 1285 950 1289
rect 954 1285 976 1289
rect 980 1285 990 1289
rect 994 1285 1008 1289
rect 1012 1285 1027 1289
rect 1031 1285 1044 1289
rect 1048 1285 1058 1289
rect 1062 1285 1065 1289
rect 1005 1206 1009 1210
rect 990 1202 994 1206
rect 998 1202 1015 1206
rect 1019 1202 1024 1206
rect 1020 1194 1024 1202
rect 990 1175 994 1190
rect 1021 1179 1051 1183
rect 974 1171 994 1175
rect 1006 1171 1041 1175
rect 885 1162 926 1166
rect 885 1149 889 1162
rect 922 1154 926 1162
rect 930 1154 947 1158
rect 951 1154 956 1158
rect 861 1145 864 1149
rect 868 1145 879 1149
rect 883 1145 889 1149
rect 952 1146 956 1154
rect 879 1137 883 1145
rect 865 1126 869 1133
rect 922 1127 926 1142
rect 974 1135 978 1171
rect 990 1167 994 1171
rect 990 1163 1009 1167
rect 1005 1154 1009 1163
rect 990 1140 994 1150
rect 1020 1140 1024 1150
rect 988 1136 996 1140
rect 1000 1136 1015 1140
rect 1019 1136 1025 1140
rect 953 1131 978 1135
rect 1037 1131 1041 1171
rect 1046 1170 1051 1179
rect 1046 1166 1101 1170
rect 1056 1158 1061 1162
rect 1065 1158 1082 1162
rect 1086 1158 1093 1162
rect 1087 1150 1091 1158
rect 1057 1131 1061 1146
rect 1096 1139 1101 1166
rect 1133 1139 1137 1312
rect 1088 1135 1112 1139
rect 1135 1135 1137 1139
rect 1037 1127 1061 1131
rect 1073 1127 1112 1131
rect 833 1122 869 1126
rect 879 1123 926 1127
rect 938 1123 978 1127
rect 833 1005 838 1122
rect 865 1115 869 1122
rect 922 1119 926 1123
rect 922 1115 941 1119
rect 879 1101 883 1111
rect 937 1106 941 1115
rect 861 1097 865 1101
rect 869 1097 879 1101
rect 883 1097 891 1101
rect 887 1092 891 1097
rect 922 1092 926 1102
rect 952 1092 956 1102
rect 974 1092 978 1123
rect 990 1119 994 1123
rect 998 1119 1015 1123
rect 1019 1119 1026 1123
rect 1020 1111 1024 1119
rect 990 1092 994 1107
rect 1037 1100 1041 1127
rect 1057 1123 1061 1127
rect 1057 1119 1076 1123
rect 1072 1110 1076 1119
rect 1021 1096 1041 1100
rect 1057 1096 1061 1106
rect 1087 1096 1091 1106
rect 1058 1092 1063 1096
rect 1067 1092 1082 1096
rect 1086 1092 1095 1096
rect 887 1088 928 1092
rect 932 1088 947 1092
rect 951 1088 958 1092
rect 974 1088 994 1092
rect 1006 1088 1032 1092
rect 1098 1088 1103 1127
rect 990 1084 994 1088
rect 1028 1084 1103 1088
rect 990 1080 1009 1084
rect 1005 1071 1009 1080
rect 990 1057 994 1067
rect 1020 1057 1024 1067
rect 988 1053 996 1057
rect 1000 1053 1015 1057
rect 1019 1053 1026 1057
rect 835 1001 838 1005
rect 885 984 890 988
rect 894 984 905 988
rect 909 984 921 988
rect 925 984 942 988
rect 946 984 967 988
rect 971 984 982 988
rect 986 984 998 988
rect 1002 984 1019 988
rect 1023 984 1035 988
rect 1039 984 1050 988
rect 1054 984 1056 988
rect 905 976 909 984
rect 947 976 951 984
rect 982 976 986 984
rect 1024 976 1028 984
rect 1050 976 1054 984
rect 891 955 895 972
rect 917 957 921 972
rect 968 957 972 972
rect 994 957 998 972
rect 1036 965 1040 972
rect 1133 966 1137 1135
rect 1150 1131 1154 1329
rect 1152 1127 1154 1131
rect 1025 961 1040 965
rect 1050 962 1056 966
rect 1135 962 1137 966
rect 794 932 796 936
rect 792 842 796 932
rect 875 951 895 955
rect 905 953 921 957
rect 933 953 972 957
rect 982 953 998 957
rect 1010 953 1025 957
rect 875 842 879 951
rect 891 936 895 951
rect 917 949 921 953
rect 917 945 936 949
rect 932 936 936 945
rect 968 936 972 953
rect 994 949 998 953
rect 1021 949 1025 953
rect 994 945 1013 949
rect 1021 945 1026 949
rect 1009 936 1013 945
rect 1036 936 1040 961
rect 1051 945 1056 949
rect 905 922 909 932
rect 917 922 921 932
rect 947 922 951 932
rect 982 922 986 932
rect 994 922 998 932
rect 1024 922 1028 932
rect 1050 922 1054 932
rect 889 918 891 922
rect 895 918 905 922
rect 909 918 923 922
rect 927 918 942 922
rect 946 918 968 922
rect 972 918 982 922
rect 986 918 1000 922
rect 1004 918 1019 922
rect 1023 918 1036 922
rect 1040 918 1050 922
rect 1054 918 1057 922
rect -43 824 -39 839
rect -17 824 -13 841
rect 22 838 131 842
rect 877 838 879 842
rect 431 835 435 838
rect 448 835 452 838
rect 775 835 779 838
rect 792 835 796 838
rect 1133 835 1137 962
rect 1150 949 1154 1127
rect 1180 1129 1184 1400
rect 1286 1278 1290 1515
rect 1304 1307 1305 1311
rect 1309 1307 1320 1311
rect 1324 1307 1336 1311
rect 1340 1307 1357 1311
rect 1361 1307 1373 1311
rect 1377 1307 1388 1311
rect 1392 1307 1394 1311
rect 1320 1299 1324 1307
rect 1362 1299 1366 1307
rect 1388 1299 1392 1307
rect 1306 1278 1310 1295
rect 1332 1280 1336 1295
rect 1374 1288 1378 1295
rect 1363 1284 1378 1288
rect 1388 1285 1394 1289
rect 1286 1274 1310 1278
rect 1320 1276 1336 1280
rect 1348 1276 1363 1280
rect 1306 1259 1310 1274
rect 1332 1272 1336 1276
rect 1359 1272 1363 1276
rect 1332 1268 1351 1272
rect 1359 1268 1364 1272
rect 1347 1259 1351 1268
rect 1374 1259 1378 1284
rect 1479 1272 1483 1313
rect 1496 1289 1500 1315
rect 1498 1285 1500 1289
rect 1389 1268 1394 1272
rect 1481 1268 1483 1272
rect 1320 1245 1324 1255
rect 1332 1245 1336 1255
rect 1362 1245 1366 1255
rect 1388 1245 1392 1255
rect 1304 1241 1306 1245
rect 1310 1241 1320 1245
rect 1324 1241 1338 1245
rect 1342 1241 1357 1245
rect 1361 1241 1374 1245
rect 1378 1241 1388 1245
rect 1392 1241 1396 1245
rect 1351 1209 1355 1213
rect 1336 1205 1340 1209
rect 1344 1205 1361 1209
rect 1365 1205 1370 1209
rect 1366 1197 1370 1205
rect 1336 1178 1340 1193
rect 1367 1182 1397 1186
rect 1320 1174 1340 1178
rect 1352 1174 1387 1178
rect 1231 1165 1272 1169
rect 1231 1152 1235 1165
rect 1268 1157 1272 1165
rect 1276 1157 1293 1161
rect 1297 1157 1302 1161
rect 1207 1148 1210 1152
rect 1214 1148 1225 1152
rect 1229 1148 1235 1152
rect 1298 1149 1302 1157
rect 1225 1140 1229 1148
rect 1211 1129 1215 1136
rect 1268 1130 1272 1145
rect 1320 1138 1324 1174
rect 1336 1170 1340 1174
rect 1336 1166 1355 1170
rect 1351 1157 1355 1166
rect 1336 1143 1340 1153
rect 1366 1143 1370 1153
rect 1334 1139 1342 1143
rect 1346 1139 1361 1143
rect 1365 1139 1371 1143
rect 1299 1134 1324 1138
rect 1383 1134 1387 1174
rect 1392 1173 1397 1182
rect 1392 1169 1447 1173
rect 1402 1161 1407 1165
rect 1411 1161 1428 1165
rect 1432 1161 1439 1165
rect 1433 1153 1437 1161
rect 1403 1134 1407 1149
rect 1442 1142 1447 1169
rect 1479 1142 1483 1268
rect 1434 1138 1458 1142
rect 1481 1138 1483 1142
rect 1383 1130 1407 1134
rect 1419 1130 1458 1134
rect 1180 1125 1215 1129
rect 1225 1126 1272 1130
rect 1284 1126 1324 1130
rect 1180 995 1184 1125
rect 1211 1118 1215 1125
rect 1268 1122 1272 1126
rect 1268 1118 1287 1122
rect 1225 1104 1229 1114
rect 1283 1109 1287 1118
rect 1207 1100 1211 1104
rect 1215 1100 1225 1104
rect 1229 1100 1237 1104
rect 1233 1095 1237 1100
rect 1268 1095 1272 1105
rect 1298 1095 1302 1105
rect 1320 1095 1324 1126
rect 1336 1122 1340 1126
rect 1344 1122 1361 1126
rect 1365 1122 1372 1126
rect 1366 1114 1370 1122
rect 1336 1095 1340 1110
rect 1383 1103 1387 1130
rect 1403 1126 1407 1130
rect 1403 1122 1422 1126
rect 1418 1113 1422 1122
rect 1367 1099 1387 1103
rect 1403 1099 1407 1109
rect 1433 1099 1437 1109
rect 1404 1095 1409 1099
rect 1413 1095 1428 1099
rect 1432 1095 1441 1099
rect 1233 1091 1274 1095
rect 1278 1091 1293 1095
rect 1297 1091 1304 1095
rect 1320 1091 1340 1095
rect 1352 1091 1378 1095
rect 1444 1091 1449 1130
rect 1336 1087 1340 1091
rect 1374 1087 1449 1091
rect 1336 1083 1355 1087
rect 1351 1074 1355 1083
rect 1336 1060 1340 1070
rect 1366 1060 1370 1070
rect 1334 1056 1342 1060
rect 1346 1056 1361 1060
rect 1365 1056 1372 1060
rect 1312 1027 1313 1031
rect 1317 1027 1328 1031
rect 1332 1027 1344 1031
rect 1348 1027 1365 1031
rect 1369 1027 1381 1031
rect 1385 1027 1396 1031
rect 1400 1027 1402 1031
rect 1328 1019 1332 1027
rect 1370 1019 1374 1027
rect 1396 1019 1400 1027
rect 1314 998 1318 1015
rect 1340 1000 1344 1015
rect 1382 1008 1386 1015
rect 1479 1009 1483 1138
rect 1496 1134 1500 1285
rect 1498 1130 1500 1134
rect 1371 1004 1386 1008
rect 1396 1005 1402 1009
rect 1481 1005 1483 1009
rect 1182 991 1184 995
rect 1293 994 1318 998
rect 1328 996 1344 1000
rect 1356 996 1371 1000
rect 1152 945 1154 949
rect 1150 835 1154 945
rect 1293 835 1297 994
rect 1314 979 1318 994
rect 1340 992 1344 996
rect 1367 992 1371 996
rect 1340 988 1359 992
rect 1367 988 1372 992
rect 1355 979 1359 988
rect 1382 979 1386 1004
rect 1397 988 1402 992
rect 1328 965 1332 975
rect 1340 965 1344 975
rect 1370 965 1374 975
rect 1396 965 1400 975
rect 1312 961 1314 965
rect 1318 961 1328 965
rect 1332 961 1346 965
rect 1350 961 1365 965
rect 1369 961 1382 965
rect 1386 961 1396 965
rect 1400 961 1404 965
rect -2 831 129 835
rect 1295 831 1297 835
rect -29 810 -25 820
rect 72 810 76 820
rect -47 806 -43 810
rect -39 806 -29 810
rect -25 806 -11 810
rect -7 806 17 810
rect 21 806 43 810
rect 47 806 67 810
rect 71 806 78 810
rect 27 779 31 806
rect 431 758 435 831
rect 448 757 452 831
rect 775 758 779 831
rect 792 757 796 831
rect 1133 757 1137 831
rect 1150 757 1154 831
rect 1479 755 1483 1005
rect 1496 992 1500 1130
rect 1498 988 1500 992
rect 1496 757 1500 988
rect -822 582 2067 584
rect -822 580 -322 582
rect -318 580 2067 582
rect -844 543 1897 545
rect -844 541 -245 543
rect -241 541 1897 543
rect -824 482 1543 484
rect -824 480 -476 482
rect -472 480 1543 482
rect -842 468 1110 470
rect -842 466 -399 468
rect -395 466 1110 468
rect 1106 446 1110 466
rect -822 377 1038 379
rect -822 375 -630 377
rect -626 375 1038 377
rect -841 358 714 360
rect -841 356 -553 358
rect -549 356 714 358
rect 710 342 714 356
rect -821 317 480 319
rect -821 315 -784 317
rect -780 315 480 317
rect -837 302 310 304
rect -837 300 -707 302
rect -703 300 306 302
rect -131 291 232 293
rect -131 289 -45 291
rect -41 289 111 291
rect 115 289 232 291
rect 133 275 140 279
rect 144 275 159 279
rect 163 275 177 279
rect 181 275 191 279
rect 195 275 199 279
rect 135 265 139 275
rect 165 265 169 275
rect 177 265 181 275
rect 150 252 154 261
rect 150 248 169 252
rect 165 244 169 248
rect 191 246 195 261
rect 140 240 153 244
rect 165 240 181 244
rect 191 242 230 246
rect 133 232 138 236
rect -796 225 -169 227
rect -796 223 -769 225
rect -765 223 -692 225
rect -688 223 -615 225
rect -611 223 -538 225
rect -534 223 -461 225
rect -457 223 -384 225
rect -380 223 -307 225
rect -303 223 -230 225
rect -226 223 -169 225
rect 165 225 169 240
rect 191 225 195 242
rect 476 222 480 315
rect -819 214 -791 218
rect -787 214 -762 218
rect -758 214 -750 218
rect -746 214 -736 218
rect -732 214 -714 218
rect -710 214 -685 218
rect -681 214 -673 218
rect -669 214 -659 218
rect -655 214 -637 218
rect -633 214 -608 218
rect -604 214 -596 218
rect -592 214 -582 218
rect -578 214 -560 218
rect -556 214 -531 218
rect -527 214 -519 218
rect -515 214 -505 218
rect -501 214 -483 218
rect -479 214 -454 218
rect -450 214 -442 218
rect -438 214 -428 218
rect -424 214 -406 218
rect -402 214 -377 218
rect -373 214 -365 218
rect -361 214 -351 218
rect -347 214 -329 218
rect -325 214 -300 218
rect -296 214 -288 218
rect -284 214 -274 218
rect -270 214 -252 218
rect -248 214 -223 218
rect -219 214 -211 218
rect -207 214 -197 218
rect -193 214 -78 218
rect -819 39 -815 214
rect -792 204 -788 214
rect -762 204 -758 214
rect -750 204 -746 214
rect -715 204 -711 214
rect -685 204 -681 214
rect -673 204 -669 214
rect -638 204 -634 214
rect -608 204 -604 214
rect -596 204 -592 214
rect -561 204 -557 214
rect -531 204 -527 214
rect -519 204 -515 214
rect -484 204 -480 214
rect -454 204 -450 214
rect -442 204 -438 214
rect -407 204 -403 214
rect -377 204 -373 214
rect -365 204 -361 214
rect -330 204 -326 214
rect -300 204 -296 214
rect -288 204 -284 214
rect -253 204 -249 214
rect -223 204 -219 214
rect -211 204 -207 214
rect -777 191 -773 200
rect -777 187 -758 191
rect -762 183 -758 187
rect -736 185 -732 200
rect -700 191 -696 200
rect -700 187 -681 191
rect -762 179 -746 183
rect -736 181 -728 185
rect -685 183 -681 187
rect -659 185 -655 200
rect -623 191 -619 200
rect -623 187 -604 191
rect -762 164 -758 179
rect -736 164 -732 181
rect -685 179 -669 183
rect -659 181 -651 185
rect -608 183 -604 187
rect -582 185 -578 200
rect -546 191 -542 200
rect -546 187 -527 191
rect -685 164 -681 179
rect -659 164 -655 181
rect -608 179 -592 183
rect -582 181 -574 185
rect -531 183 -527 187
rect -505 185 -501 200
rect -469 191 -465 200
rect -469 187 -450 191
rect -608 164 -604 179
rect -582 164 -578 181
rect -531 179 -515 183
rect -505 181 -497 185
rect -454 183 -450 187
rect -428 185 -424 200
rect -392 191 -388 200
rect -392 187 -373 191
rect -531 164 -527 179
rect -505 164 -501 181
rect -454 179 -438 183
rect -428 181 -420 185
rect -377 183 -373 187
rect -351 185 -347 200
rect -315 191 -311 200
rect -315 187 -296 191
rect -454 164 -450 179
rect -428 164 -424 181
rect -377 179 -361 183
rect -351 181 -343 185
rect -300 183 -296 187
rect -274 185 -270 200
rect -238 191 -234 200
rect -238 187 -219 191
rect -377 164 -373 179
rect -351 164 -347 181
rect -300 179 -284 183
rect -274 181 -266 185
rect -223 183 -219 187
rect -197 185 -193 200
rect -82 203 -78 214
rect 135 213 139 221
rect 177 213 181 221
rect 1034 219 1038 375
rect 1539 219 1543 480
rect 133 209 140 213
rect 144 209 161 213
rect 165 209 177 213
rect 181 209 192 213
rect 196 209 197 213
rect 238 210 2104 212
rect 238 208 441 210
rect 445 208 800 210
rect 804 208 999 210
rect 1003 208 1305 210
rect 1309 208 1504 210
rect 1508 208 1829 210
rect 1833 208 2028 210
rect 2032 208 2104 210
rect -82 199 -71 203
rect -67 199 -57 203
rect -53 199 -51 203
rect 135 199 142 203
rect 146 199 161 203
rect 165 199 179 203
rect 183 199 193 203
rect 197 199 288 203
rect 292 199 313 203
rect 317 199 325 203
rect 329 199 339 203
rect 343 199 458 203
rect 462 199 483 203
rect 487 199 495 203
rect 499 199 509 203
rect 513 199 846 203
rect 850 199 871 203
rect 875 199 883 203
rect 887 199 897 203
rect 901 199 1016 203
rect 1020 199 1041 203
rect 1045 199 1053 203
rect 1057 199 1067 203
rect 1071 199 1351 203
rect 1355 199 1376 203
rect 1380 199 1388 203
rect 1392 199 1402 203
rect 1406 199 1521 203
rect 1525 199 1546 203
rect 1550 199 1558 203
rect 1562 199 1572 203
rect 1576 199 1875 203
rect 1879 199 1900 203
rect 1904 199 1912 203
rect 1916 199 1926 203
rect 1930 199 2045 203
rect 2049 199 2070 203
rect 2074 199 2082 203
rect 2086 199 2096 203
rect 2100 199 2104 203
rect -71 189 -67 199
rect 137 189 141 199
rect 167 189 171 199
rect 179 189 183 199
rect 283 189 287 199
rect 313 189 317 199
rect 325 189 329 199
rect 453 189 457 199
rect 483 189 487 199
rect 495 189 499 199
rect 841 189 845 199
rect 871 189 875 199
rect 883 189 887 199
rect 1011 189 1015 199
rect 1041 189 1045 199
rect 1053 189 1057 199
rect 1346 189 1350 199
rect 1376 189 1380 199
rect 1388 189 1392 199
rect 1516 189 1520 199
rect 1546 189 1550 199
rect 1558 189 1562 199
rect 1870 189 1874 199
rect 1900 189 1904 199
rect 1912 189 1916 199
rect 2040 189 2044 199
rect 2070 189 2074 199
rect 2082 189 2086 199
rect -300 164 -296 179
rect -274 164 -270 181
rect -223 179 -207 183
rect -197 181 -189 185
rect -223 164 -219 179
rect -197 164 -193 181
rect -57 170 -53 185
rect 152 176 156 185
rect 152 172 171 176
rect -131 164 -67 168
rect -57 166 61 170
rect 167 168 171 172
rect 193 170 197 185
rect 298 176 302 185
rect 298 172 317 176
rect -792 152 -788 160
rect -750 152 -746 160
rect -715 152 -711 160
rect -673 152 -669 160
rect -638 152 -634 160
rect -596 152 -592 160
rect -561 152 -557 160
rect -519 152 -515 160
rect -484 152 -480 160
rect -442 152 -438 160
rect -407 152 -403 160
rect -365 152 -361 160
rect -330 152 -326 160
rect -288 152 -284 160
rect -253 152 -249 160
rect -211 152 -207 160
rect -796 148 -787 152
rect -783 148 -766 152
rect -762 148 -750 152
rect -746 148 -735 152
rect -731 148 -710 152
rect -706 148 -689 152
rect -685 148 -673 152
rect -669 148 -658 152
rect -654 148 -633 152
rect -629 148 -612 152
rect -608 148 -596 152
rect -592 148 -581 152
rect -577 148 -556 152
rect -552 148 -535 152
rect -531 148 -519 152
rect -515 148 -504 152
rect -500 148 -479 152
rect -475 148 -458 152
rect -454 148 -442 152
rect -438 148 -427 152
rect -423 148 -402 152
rect -398 148 -381 152
rect -377 148 -365 152
rect -361 148 -350 152
rect -346 148 -325 152
rect -321 148 -304 152
rect -300 148 -288 152
rect -284 148 -273 152
rect -269 148 -248 152
rect -244 148 -227 152
rect -223 148 -211 152
rect -207 148 -196 152
rect -192 148 -172 152
rect -91 128 -87 164
rect -57 149 -53 166
rect 94 164 155 168
rect 167 164 183 168
rect 193 166 230 170
rect 313 168 317 172
rect 339 170 343 185
rect 468 176 472 185
rect 468 172 487 176
rect 94 145 98 164
rect -71 137 -67 145
rect 56 141 98 145
rect 125 156 140 160
rect -72 133 -71 137
rect -67 133 -56 137
rect -52 133 -49 137
rect -91 126 34 128
rect 56 128 60 141
rect 38 126 60 128
rect -91 124 60 126
rect -74 115 -71 119
rect -67 115 -57 119
rect -53 115 -51 119
rect -71 105 -67 115
rect 125 113 129 156
rect 167 149 171 164
rect 193 149 197 166
rect 313 164 329 168
rect 339 166 349 170
rect 483 168 487 172
rect 509 170 513 185
rect 856 176 860 185
rect 856 172 875 176
rect 313 149 317 164
rect 339 149 343 166
rect 483 164 499 168
rect 509 166 519 170
rect 871 168 875 172
rect 897 170 901 185
rect 1026 176 1030 185
rect 1026 172 1045 176
rect 483 149 487 164
rect 509 149 513 166
rect 871 164 887 168
rect 897 166 907 170
rect 1041 168 1045 172
rect 1067 170 1071 185
rect 1361 176 1365 185
rect 1361 172 1380 176
rect 871 149 875 164
rect 897 149 901 166
rect 1041 164 1057 168
rect 1067 166 1077 170
rect 1376 168 1380 172
rect 1402 170 1406 185
rect 1531 176 1535 185
rect 1531 172 1550 176
rect 1041 149 1045 164
rect 1067 149 1071 166
rect 1376 164 1392 168
rect 1402 166 1412 170
rect 1546 168 1550 172
rect 1572 170 1576 185
rect 1885 176 1889 185
rect 1885 172 1904 176
rect 1376 149 1380 164
rect 1402 149 1406 166
rect 1546 164 1562 168
rect 1572 166 1582 170
rect 1900 168 1904 172
rect 1926 170 1930 185
rect 2055 176 2059 185
rect 2055 172 2074 176
rect 1546 149 1550 164
rect 1572 149 1576 166
rect 1900 164 1916 168
rect 1926 166 1936 170
rect 2070 168 2074 172
rect 2096 170 2100 185
rect 1900 149 1904 164
rect 1926 149 1930 166
rect 2070 164 2086 168
rect 2096 166 2106 170
rect 2070 149 2074 164
rect 2096 149 2100 166
rect 137 137 141 145
rect 179 137 183 145
rect 283 137 287 145
rect 325 137 329 145
rect 453 137 457 145
rect 495 137 499 145
rect 841 137 845 145
rect 883 137 887 145
rect 1011 137 1015 145
rect 1053 137 1057 145
rect 1346 137 1350 145
rect 1388 137 1392 145
rect 1516 137 1520 145
rect 1558 137 1562 145
rect 1870 137 1874 145
rect 1912 137 1916 145
rect 2040 137 2044 145
rect 2082 137 2086 145
rect 135 133 142 137
rect 146 133 163 137
rect 167 133 179 137
rect 183 133 194 137
rect 198 133 199 137
rect 234 133 284 137
rect 288 133 312 137
rect 316 133 325 137
rect 329 133 340 137
rect 344 133 454 137
rect 458 133 482 137
rect 486 133 495 137
rect 499 133 510 137
rect 514 133 842 137
rect 846 133 870 137
rect 874 133 883 137
rect 887 133 898 137
rect 902 133 1012 137
rect 1016 133 1040 137
rect 1044 133 1053 137
rect 1057 133 1068 137
rect 1072 133 1347 137
rect 1351 133 1375 137
rect 1379 133 1388 137
rect 1392 133 1403 137
rect 1407 133 1517 137
rect 1521 133 1545 137
rect 1549 133 1558 137
rect 1562 133 1573 137
rect 1577 133 1871 137
rect 1875 133 1899 137
rect 1903 133 1912 137
rect 1916 133 1927 137
rect 1931 133 2041 137
rect 2045 133 2069 137
rect 2073 133 2082 137
rect 2086 133 2097 137
rect 2101 133 2104 137
rect 137 123 144 127
rect 148 123 163 127
rect 167 123 181 127
rect 185 123 195 127
rect 199 123 268 127
rect 58 109 129 113
rect 139 113 143 123
rect 169 113 173 123
rect 181 113 185 123
rect -57 86 -53 101
rect 58 86 62 109
rect 154 100 158 109
rect 137 96 146 100
rect 154 96 173 100
rect 142 92 146 96
rect 169 92 173 96
rect 195 94 199 109
rect 142 88 157 92
rect 169 88 185 92
rect 195 90 250 94
rect -57 84 62 86
rect -131 80 -67 84
rect -57 82 58 84
rect -91 45 -87 80
rect -57 65 -53 82
rect 75 80 142 84
rect -71 53 -67 61
rect -72 49 -71 53
rect -67 49 -56 53
rect -52 49 -49 53
rect 75 45 79 80
rect 169 73 173 88
rect 195 73 199 90
rect 139 61 143 69
rect 181 61 185 69
rect 246 62 250 90
rect 264 89 268 123
rect 345 96 2211 98
rect 345 94 548 96
rect 552 94 907 96
rect 911 94 1106 96
rect 1110 94 1412 96
rect 1416 94 1611 96
rect 1615 94 1936 96
rect 1940 94 2135 96
rect 2139 94 2211 96
rect 264 85 273 89
rect 277 85 292 89
rect 296 85 310 89
rect 314 85 324 89
rect 328 85 395 89
rect 399 85 420 89
rect 424 85 432 89
rect 436 85 446 89
rect 450 85 565 89
rect 569 85 590 89
rect 594 85 602 89
rect 606 85 616 89
rect 620 85 953 89
rect 957 85 978 89
rect 982 85 990 89
rect 994 85 1004 89
rect 1008 85 1123 89
rect 1127 85 1148 89
rect 1152 85 1160 89
rect 1164 85 1174 89
rect 1178 85 1458 89
rect 1462 85 1483 89
rect 1487 85 1495 89
rect 1499 85 1509 89
rect 1513 85 1628 89
rect 1632 85 1653 89
rect 1657 85 1665 89
rect 1669 85 1679 89
rect 1683 85 1982 89
rect 1986 85 2007 89
rect 2011 85 2019 89
rect 2023 85 2033 89
rect 2037 85 2152 89
rect 2156 85 2177 89
rect 2181 85 2189 89
rect 2193 85 2203 89
rect 2207 85 2255 89
rect 268 75 272 85
rect 310 75 314 85
rect 390 75 394 85
rect 420 75 424 85
rect 432 75 436 85
rect 560 75 564 85
rect 590 75 594 85
rect 602 75 606 85
rect 948 75 952 85
rect 978 75 982 85
rect 990 75 994 85
rect 1118 75 1122 85
rect 1148 75 1152 85
rect 1160 75 1164 85
rect 1453 75 1457 85
rect 1483 75 1487 85
rect 1495 75 1499 85
rect 1623 75 1627 85
rect 1653 75 1657 85
rect 1665 75 1669 85
rect 1977 75 1981 85
rect 2007 75 2011 85
rect 2019 75 2023 85
rect 2147 75 2151 85
rect 2177 75 2181 85
rect 2189 75 2193 85
rect 137 57 144 61
rect 148 57 165 61
rect 169 57 181 61
rect 185 57 196 61
rect 200 57 201 61
rect 246 58 287 62
rect 298 54 302 71
rect 324 56 328 71
rect 405 62 409 71
rect 405 58 424 62
rect 139 47 146 51
rect 150 47 165 51
rect 169 47 183 51
rect 187 47 197 51
rect 201 47 203 51
rect 282 50 314 54
rect 324 52 330 56
rect 420 54 424 58
rect 446 56 450 71
rect 575 62 579 71
rect 575 58 594 62
rect -91 41 79 45
rect -819 35 -612 39
rect -608 35 -593 39
rect -589 35 -575 39
rect -571 35 -561 39
rect -557 35 -535 39
rect -531 35 -516 39
rect -512 35 -498 39
rect -494 35 -484 39
rect -480 35 -458 39
rect -454 35 -439 39
rect -435 35 -421 39
rect -417 35 -407 39
rect -403 35 -381 39
rect -377 35 -362 39
rect -358 35 -344 39
rect -340 35 -330 39
rect -326 35 -322 39
rect 141 37 145 47
rect 171 37 175 47
rect -617 25 -613 35
rect -587 25 -583 35
rect -575 25 -571 35
rect -540 25 -536 35
rect -510 25 -506 35
rect -498 25 -494 35
rect -463 25 -459 35
rect -433 25 -429 35
rect -421 25 -417 35
rect -386 25 -382 35
rect -356 25 -352 35
rect -344 25 -340 35
rect 183 37 187 47
rect 228 42 271 46
rect -602 12 -598 21
rect -602 8 -583 12
rect -587 4 -583 8
rect -561 6 -557 21
rect -525 12 -521 21
rect -525 8 -506 12
rect -587 0 -571 4
rect -561 2 -555 6
rect -510 4 -506 8
rect -484 6 -480 21
rect -448 12 -444 21
rect -448 8 -429 12
rect -587 -15 -583 0
rect -561 -15 -557 2
rect -510 0 -494 4
rect -484 2 -478 6
rect -433 4 -429 8
rect -407 6 -403 21
rect -371 12 -367 21
rect -371 8 -352 12
rect -510 -15 -506 0
rect -484 -15 -480 2
rect -433 0 -417 4
rect -407 2 -401 6
rect -356 4 -352 8
rect -330 6 -326 21
rect 156 24 160 33
rect 156 20 175 24
rect 171 16 175 20
rect 197 18 201 33
rect 228 18 232 42
rect 282 35 286 50
rect 324 35 328 52
rect 420 50 436 54
rect 446 52 456 56
rect 590 54 594 58
rect 616 56 620 71
rect 963 62 967 71
rect 963 58 982 62
rect 420 35 424 50
rect 446 35 450 52
rect 590 50 606 54
rect 616 52 626 56
rect 978 54 982 58
rect 1004 56 1008 71
rect 1133 62 1137 71
rect 1133 58 1152 62
rect 590 35 594 50
rect 616 35 620 52
rect 978 50 994 54
rect 1004 52 1014 56
rect 1148 54 1152 58
rect 1174 56 1178 71
rect 1468 62 1472 71
rect 1468 58 1487 62
rect 978 35 982 50
rect 1004 35 1008 52
rect 1148 50 1164 54
rect 1174 52 1184 56
rect 1483 54 1487 58
rect 1509 56 1513 71
rect 1638 62 1642 71
rect 1638 58 1657 62
rect 1148 35 1152 50
rect 1174 35 1178 52
rect 1483 50 1499 54
rect 1509 52 1519 56
rect 1653 54 1657 58
rect 1679 56 1683 71
rect 1992 62 1996 71
rect 1992 58 2011 62
rect 1483 35 1487 50
rect 1509 35 1513 52
rect 1653 50 1669 54
rect 1679 52 1689 56
rect 2007 54 2011 58
rect 2033 56 2037 71
rect 2162 62 2166 71
rect 2162 58 2181 62
rect 1653 35 1657 50
rect 1679 35 1683 52
rect 2007 50 2023 54
rect 2033 52 2043 56
rect 2177 54 2181 58
rect 2203 56 2207 71
rect 2007 35 2011 50
rect 2033 35 2037 52
rect 2177 50 2193 54
rect 2203 52 2213 56
rect 2177 35 2181 50
rect 2203 35 2207 52
rect 268 23 272 31
rect 298 23 302 31
rect 310 23 314 31
rect 390 23 394 31
rect 432 23 436 31
rect 560 23 564 31
rect 602 23 606 31
rect 948 23 952 31
rect 990 23 994 31
rect 1118 23 1122 31
rect 1160 23 1164 31
rect 1453 23 1457 31
rect 1495 23 1499 31
rect 1623 23 1627 31
rect 1665 23 1669 31
rect 1977 23 1981 31
rect 2019 23 2023 31
rect 2147 23 2151 31
rect 2189 23 2193 31
rect 268 19 273 23
rect 277 19 294 23
rect 298 19 310 23
rect 314 19 325 23
rect 329 19 391 23
rect 395 19 419 23
rect 423 19 432 23
rect 436 19 447 23
rect 451 19 561 23
rect 565 19 589 23
rect 593 19 602 23
rect 606 19 617 23
rect 621 19 949 23
rect 953 19 977 23
rect 981 19 990 23
rect 994 19 1005 23
rect 1009 19 1119 23
rect 1123 19 1147 23
rect 1151 19 1160 23
rect 1164 19 1175 23
rect 1179 19 1454 23
rect 1458 19 1482 23
rect 1486 19 1495 23
rect 1499 19 1510 23
rect 1514 19 1624 23
rect 1628 19 1652 23
rect 1656 19 1665 23
rect 1669 19 1680 23
rect 1684 19 1978 23
rect 1982 19 2006 23
rect 2010 19 2019 23
rect 2023 19 2034 23
rect 2038 19 2148 23
rect 2152 19 2176 23
rect 2180 19 2189 23
rect 2193 19 2204 23
rect 2208 19 2211 23
rect 146 12 159 16
rect 171 12 187 16
rect 197 14 232 18
rect 62 6 144 8
rect -433 -15 -429 0
rect -407 -15 -403 2
rect -356 0 -340 4
rect -330 2 -324 6
rect 58 4 144 6
rect -356 -15 -352 0
rect -330 -15 -326 2
rect 171 -3 175 12
rect 197 -3 201 14
rect 141 -15 145 -7
rect 183 -15 187 -7
rect 139 -19 146 -15
rect 150 -19 167 -15
rect 171 -19 183 -15
rect 187 -19 198 -15
rect 202 -19 203 -15
rect -617 -27 -613 -19
rect -575 -27 -571 -19
rect -540 -27 -536 -19
rect -498 -27 -494 -19
rect -463 -27 -459 -19
rect -421 -27 -417 -19
rect -386 -27 -382 -19
rect -344 -27 -340 -19
rect -618 -31 -612 -27
rect -608 -31 -591 -27
rect -587 -31 -575 -27
rect -571 -31 -560 -27
rect -556 -31 -535 -27
rect -531 -31 -514 -27
rect -510 -31 -498 -27
rect -494 -31 -483 -27
rect -479 -31 -458 -27
rect -454 -31 -437 -27
rect -433 -31 -421 -27
rect -417 -31 -406 -27
rect -402 -31 -381 -27
rect -377 -31 -360 -27
rect -356 -31 -344 -27
rect -340 -31 -329 -27
rect -325 -31 -322 -27
rect -131 -28 -82 -26
rect -78 -28 216 -26
rect 220 -28 225 -26
rect -131 -30 225 -28
rect 2251 -47 2255 85
rect 395 -49 492 -47
rect 395 -51 455 -49
rect 459 -51 492 -49
rect 496 -51 511 -47
rect 515 -49 1005 -47
rect 515 -51 968 -49
rect 487 -61 491 -51
rect 517 -61 521 -51
rect 502 -74 506 -65
rect 502 -78 521 -74
rect 408 -82 483 -78
rect 517 -82 521 -78
rect 572 -82 576 -51
rect 972 -51 1005 -49
rect 1009 -51 1024 -47
rect 1028 -49 1511 -47
rect 1028 -51 1474 -49
rect 1000 -61 1004 -51
rect 1030 -61 1034 -51
rect 1015 -74 1019 -65
rect 1015 -78 1034 -74
rect 921 -82 996 -78
rect 1030 -82 1034 -78
rect 1085 -82 1089 -51
rect 1478 -51 1511 -49
rect 1515 -51 1530 -47
rect 1534 -49 2035 -47
rect 1534 -51 1998 -49
rect 1506 -61 1510 -51
rect 1536 -61 1540 -51
rect 1521 -74 1525 -65
rect 1521 -78 1540 -74
rect 1427 -82 1502 -78
rect 1536 -82 1540 -78
rect 1591 -82 1595 -51
rect 2002 -51 2035 -49
rect 2039 -51 2054 -47
rect 2058 -51 2706 -47
rect 2030 -61 2034 -51
rect 2060 -61 2064 -51
rect 2045 -74 2049 -65
rect 2045 -78 2064 -74
rect 1951 -82 2026 -78
rect 2060 -82 2064 -78
rect 2115 -82 2119 -51
rect 408 -121 413 -82
rect 479 -86 505 -82
rect 517 -86 537 -82
rect 553 -86 560 -82
rect 564 -86 579 -82
rect 583 -86 593 -82
rect 416 -90 425 -86
rect 429 -90 444 -86
rect 448 -90 453 -86
rect 420 -100 424 -90
rect 450 -100 454 -90
rect 470 -94 490 -90
rect 435 -113 439 -104
rect 435 -117 454 -113
rect 450 -121 454 -117
rect 470 -121 474 -94
rect 517 -101 521 -86
rect 487 -113 491 -105
rect 485 -117 492 -113
rect 496 -117 513 -113
rect 517 -117 521 -113
rect 533 -117 537 -86
rect 555 -96 559 -86
rect 585 -96 589 -86
rect 570 -109 574 -100
rect 570 -113 589 -109
rect 585 -117 589 -113
rect 533 -121 573 -117
rect 585 -119 640 -117
rect 585 -121 636 -119
rect 399 -125 438 -121
rect 450 -125 474 -121
rect 384 -133 423 -129
rect 384 -213 388 -133
rect 410 -160 415 -133
rect 450 -140 454 -125
rect 420 -152 424 -144
rect 418 -156 425 -152
rect 429 -156 446 -152
rect 450 -156 455 -152
rect 410 -164 465 -160
rect 460 -173 465 -164
rect 470 -165 474 -125
rect 533 -129 558 -125
rect 486 -134 492 -130
rect 496 -134 511 -130
rect 515 -134 523 -130
rect 487 -144 491 -134
rect 517 -144 521 -134
rect 502 -157 506 -148
rect 502 -161 521 -157
rect 517 -165 521 -161
rect 533 -165 537 -129
rect 585 -136 589 -121
rect 921 -121 926 -82
rect 992 -86 1018 -82
rect 1030 -86 1050 -82
rect 1066 -86 1073 -82
rect 1077 -86 1092 -82
rect 1096 -86 1106 -82
rect 929 -90 938 -86
rect 942 -90 957 -86
rect 961 -90 966 -86
rect 933 -100 937 -90
rect 963 -100 967 -90
rect 983 -94 1003 -90
rect 948 -113 952 -104
rect 948 -117 967 -113
rect 963 -121 967 -117
rect 983 -121 987 -94
rect 1030 -101 1034 -86
rect 1000 -113 1004 -105
rect 998 -117 1005 -113
rect 1009 -117 1026 -113
rect 1030 -117 1034 -113
rect 1046 -117 1050 -86
rect 1068 -96 1072 -86
rect 1098 -96 1102 -86
rect 1083 -109 1087 -100
rect 1083 -113 1102 -109
rect 1098 -117 1102 -113
rect 1046 -121 1086 -117
rect 1098 -119 1163 -117
rect 1098 -121 1159 -119
rect 912 -125 951 -121
rect 963 -125 987 -121
rect 912 -133 936 -129
rect 555 -148 559 -140
rect 555 -152 560 -148
rect 564 -152 581 -148
rect 585 -152 589 -148
rect 923 -160 928 -133
rect 963 -140 967 -125
rect 933 -152 937 -144
rect 931 -156 938 -152
rect 942 -156 959 -152
rect 963 -156 968 -152
rect 923 -164 978 -160
rect 470 -169 505 -165
rect 517 -169 537 -165
rect 460 -177 490 -173
rect 517 -184 521 -169
rect 973 -173 978 -164
rect 983 -165 987 -125
rect 1046 -129 1071 -125
rect 999 -134 1005 -130
rect 1009 -134 1024 -130
rect 1028 -134 1036 -130
rect 1000 -144 1004 -134
rect 1030 -144 1034 -134
rect 1015 -157 1019 -148
rect 1015 -161 1034 -157
rect 1030 -165 1034 -161
rect 1046 -165 1050 -129
rect 1098 -136 1102 -121
rect 1427 -121 1432 -82
rect 1498 -86 1524 -82
rect 1536 -86 1556 -82
rect 1572 -86 1579 -82
rect 1583 -86 1598 -82
rect 1602 -86 1612 -82
rect 1435 -90 1444 -86
rect 1448 -90 1463 -86
rect 1467 -90 1472 -86
rect 1439 -100 1443 -90
rect 1469 -100 1473 -90
rect 1489 -94 1509 -90
rect 1454 -113 1458 -104
rect 1454 -117 1473 -113
rect 1469 -121 1473 -117
rect 1489 -121 1493 -94
rect 1536 -101 1540 -86
rect 1506 -113 1510 -105
rect 1504 -117 1511 -113
rect 1515 -117 1532 -113
rect 1536 -117 1540 -113
rect 1552 -117 1556 -86
rect 1574 -96 1578 -86
rect 1604 -96 1608 -86
rect 1589 -109 1593 -100
rect 1589 -113 1608 -109
rect 1604 -117 1608 -113
rect 1552 -121 1592 -117
rect 1604 -119 1686 -117
rect 1604 -121 1682 -119
rect 1418 -125 1457 -121
rect 1469 -125 1493 -121
rect 1418 -133 1442 -129
rect 1068 -148 1072 -140
rect 1068 -152 1073 -148
rect 1077 -152 1094 -148
rect 1098 -152 1102 -148
rect 1429 -160 1434 -133
rect 1469 -140 1473 -125
rect 1439 -152 1443 -144
rect 1437 -156 1444 -152
rect 1448 -156 1465 -152
rect 1469 -156 1474 -152
rect 1429 -164 1484 -160
rect 983 -169 1018 -165
rect 1030 -169 1050 -165
rect 973 -177 1003 -173
rect 1030 -184 1034 -169
rect 1479 -173 1484 -164
rect 1489 -165 1493 -125
rect 1552 -129 1577 -125
rect 1505 -134 1511 -130
rect 1515 -134 1530 -130
rect 1534 -134 1542 -130
rect 1506 -144 1510 -134
rect 1536 -144 1540 -134
rect 1521 -157 1525 -148
rect 1521 -161 1540 -157
rect 1536 -165 1540 -161
rect 1552 -165 1556 -129
rect 1604 -136 1608 -121
rect 1951 -121 1956 -82
rect 2022 -86 2048 -82
rect 2060 -86 2080 -82
rect 2096 -86 2103 -82
rect 2107 -86 2122 -82
rect 2126 -86 2136 -82
rect 1959 -90 1968 -86
rect 1972 -90 1987 -86
rect 1991 -90 1996 -86
rect 1963 -100 1967 -90
rect 1993 -100 1997 -90
rect 2013 -94 2033 -90
rect 1978 -113 1982 -104
rect 1978 -117 1997 -113
rect 1993 -121 1997 -117
rect 2013 -121 2017 -94
rect 2060 -101 2064 -86
rect 2030 -113 2034 -105
rect 2028 -117 2035 -113
rect 2039 -117 2056 -113
rect 2060 -117 2064 -113
rect 2076 -117 2080 -86
rect 2098 -96 2102 -86
rect 2128 -96 2132 -86
rect 2113 -109 2117 -100
rect 2113 -113 2132 -109
rect 2128 -117 2132 -113
rect 2076 -121 2116 -117
rect 2128 -119 2209 -117
rect 2128 -121 2205 -119
rect 1942 -125 1981 -121
rect 1993 -125 2017 -121
rect 1942 -133 1966 -129
rect 1574 -148 1578 -140
rect 1574 -152 1579 -148
rect 1583 -152 1600 -148
rect 1604 -152 1608 -148
rect 1953 -160 1958 -133
rect 1993 -140 1997 -125
rect 1963 -152 1967 -144
rect 1961 -156 1968 -152
rect 1972 -156 1989 -152
rect 1993 -156 1998 -152
rect 1953 -164 2008 -160
rect 1489 -169 1524 -165
rect 1536 -169 1556 -165
rect 1479 -177 1509 -173
rect 1536 -184 1540 -169
rect 2003 -173 2008 -164
rect 2013 -165 2017 -125
rect 2076 -129 2101 -125
rect 2029 -134 2035 -130
rect 2039 -134 2054 -130
rect 2058 -134 2066 -130
rect 2030 -144 2034 -134
rect 2060 -144 2064 -134
rect 2045 -157 2049 -148
rect 2045 -161 2064 -157
rect 2060 -165 2064 -161
rect 2076 -165 2080 -129
rect 2128 -136 2132 -121
rect 2098 -148 2102 -140
rect 2098 -152 2103 -148
rect 2107 -152 2124 -148
rect 2128 -152 2132 -148
rect 2013 -169 2048 -165
rect 2060 -169 2080 -165
rect 2003 -177 2033 -173
rect 2060 -184 2064 -169
rect 395 -198 465 -196
rect 487 -196 491 -188
rect 469 -198 492 -196
rect 395 -200 492 -198
rect 496 -200 513 -196
rect 517 -198 525 -196
rect 529 -198 549 -196
rect 553 -198 978 -196
rect 1000 -196 1004 -188
rect 982 -198 1005 -196
rect 517 -200 590 -198
rect 594 -200 1005 -198
rect 1009 -200 1026 -196
rect 1030 -198 1038 -196
rect 1042 -198 1062 -196
rect 1066 -198 1484 -196
rect 1506 -196 1510 -188
rect 1488 -198 1511 -196
rect 1030 -200 1511 -198
rect 1515 -200 1532 -196
rect 1536 -198 1544 -196
rect 1548 -198 1568 -196
rect 1572 -198 2008 -196
rect 2030 -196 2034 -188
rect 2012 -198 2035 -196
rect 1536 -200 2035 -198
rect 2039 -200 2056 -196
rect 2060 -198 2068 -196
rect 2072 -198 2092 -196
rect 2096 -198 2282 -196
rect 2060 -200 2282 -198
rect 381 -215 906 -213
rect 910 -215 1412 -213
rect 1416 -215 1936 -213
rect 1940 -215 2282 -213
rect 381 -217 2282 -215
rect 462 -392 466 -217
rect 2702 -231 2706 -51
rect 614 -233 759 -231
rect 614 -235 722 -233
rect 726 -235 759 -233
rect 763 -235 778 -231
rect 782 -233 994 -231
rect 782 -235 957 -233
rect 754 -245 758 -235
rect 784 -245 788 -235
rect 769 -258 773 -249
rect 769 -262 788 -258
rect 675 -266 750 -262
rect 784 -266 788 -262
rect 839 -266 843 -235
rect 961 -235 994 -233
rect 998 -235 1013 -231
rect 1017 -233 1282 -231
rect 1017 -235 1113 -233
rect 989 -245 993 -235
rect 1019 -245 1023 -235
rect 1004 -258 1008 -249
rect 1004 -262 1023 -258
rect 910 -266 985 -262
rect 1019 -266 1023 -262
rect 1074 -266 1078 -235
rect 1117 -235 1245 -233
rect 1249 -235 1282 -233
rect 1286 -235 1301 -231
rect 1305 -233 1517 -231
rect 1305 -235 1480 -233
rect 1277 -245 1281 -235
rect 1307 -245 1311 -235
rect 1292 -258 1296 -249
rect 1292 -262 1311 -258
rect 1198 -266 1273 -262
rect 1307 -266 1311 -262
rect 1362 -266 1366 -235
rect 1484 -235 1517 -233
rect 1521 -235 1536 -231
rect 1540 -233 1805 -231
rect 1540 -235 1636 -233
rect 1512 -245 1516 -235
rect 1542 -245 1546 -235
rect 1527 -258 1531 -249
rect 1527 -262 1546 -258
rect 1433 -266 1508 -262
rect 1542 -266 1546 -262
rect 1597 -266 1601 -235
rect 1640 -235 1768 -233
rect 1772 -235 1805 -233
rect 1809 -235 1824 -231
rect 1828 -233 2040 -231
rect 1828 -235 2003 -233
rect 1800 -245 1804 -235
rect 1830 -245 1834 -235
rect 1815 -258 1819 -249
rect 1815 -262 1834 -258
rect 1721 -266 1796 -262
rect 1830 -266 1834 -262
rect 1885 -266 1889 -235
rect 2007 -235 2040 -233
rect 2044 -235 2059 -231
rect 2063 -233 2328 -231
rect 2063 -235 2159 -233
rect 2035 -245 2039 -235
rect 2065 -245 2069 -235
rect 2050 -258 2054 -249
rect 2050 -262 2069 -258
rect 1956 -266 2031 -262
rect 2065 -266 2069 -262
rect 2120 -266 2124 -235
rect 2163 -235 2291 -233
rect 2295 -235 2328 -233
rect 2332 -235 2347 -231
rect 2351 -233 2563 -231
rect 2351 -235 2526 -233
rect 2323 -245 2327 -235
rect 2353 -245 2357 -235
rect 2338 -258 2342 -249
rect 2338 -262 2357 -258
rect 2244 -266 2319 -262
rect 2353 -266 2357 -262
rect 2408 -266 2412 -235
rect 2530 -235 2563 -233
rect 2567 -235 2582 -231
rect 2586 -233 2706 -231
rect 2586 -235 2682 -233
rect 2558 -245 2562 -235
rect 2588 -245 2592 -235
rect 2573 -258 2577 -249
rect 2573 -262 2592 -258
rect 2479 -266 2554 -262
rect 2588 -266 2592 -262
rect 2643 -266 2647 -235
rect 2686 -235 2706 -233
rect 640 -307 662 -305
rect 675 -305 680 -266
rect 746 -270 772 -266
rect 784 -270 804 -266
rect 820 -270 827 -266
rect 831 -270 846 -266
rect 850 -270 860 -266
rect 683 -274 692 -270
rect 696 -274 711 -270
rect 715 -274 720 -270
rect 687 -284 691 -274
rect 717 -284 721 -274
rect 737 -278 757 -274
rect 702 -297 706 -288
rect 702 -301 721 -297
rect 717 -305 721 -301
rect 737 -305 741 -278
rect 784 -285 788 -270
rect 754 -297 758 -289
rect 752 -301 759 -297
rect 763 -301 780 -297
rect 784 -301 788 -297
rect 800 -301 804 -270
rect 822 -280 826 -270
rect 852 -280 856 -270
rect 837 -293 841 -284
rect 837 -297 856 -293
rect 852 -301 856 -297
rect 910 -301 915 -266
rect 981 -270 1007 -266
rect 1019 -270 1039 -266
rect 1055 -270 1062 -266
rect 1066 -270 1081 -266
rect 1085 -270 1095 -266
rect 918 -274 927 -270
rect 931 -274 946 -270
rect 950 -274 955 -270
rect 922 -284 926 -274
rect 952 -284 956 -274
rect 972 -278 992 -274
rect 937 -297 941 -288
rect 937 -301 956 -297
rect 800 -305 840 -301
rect 852 -303 915 -301
rect 852 -305 881 -303
rect 666 -307 705 -305
rect 636 -309 705 -307
rect 717 -309 741 -305
rect 626 -315 628 -313
rect 632 -315 690 -313
rect 626 -317 662 -315
rect 666 -317 690 -315
rect 677 -344 682 -317
rect 717 -324 721 -309
rect 687 -336 691 -328
rect 685 -340 692 -336
rect 696 -340 713 -336
rect 717 -340 722 -336
rect 677 -348 732 -344
rect 727 -357 732 -348
rect 737 -349 741 -309
rect 800 -313 825 -309
rect 753 -318 759 -314
rect 763 -318 778 -314
rect 782 -318 790 -314
rect 754 -328 758 -318
rect 784 -328 788 -318
rect 769 -341 773 -332
rect 769 -345 788 -341
rect 784 -349 788 -345
rect 800 -349 804 -313
rect 852 -320 856 -305
rect 885 -305 915 -303
rect 952 -305 956 -301
rect 972 -305 976 -278
rect 1019 -285 1023 -270
rect 989 -297 993 -289
rect 987 -301 994 -297
rect 998 -301 1015 -297
rect 1019 -301 1023 -297
rect 1035 -301 1039 -270
rect 1057 -280 1061 -270
rect 1087 -280 1091 -270
rect 1072 -293 1076 -284
rect 1072 -297 1091 -293
rect 1087 -301 1091 -297
rect 1035 -305 1075 -301
rect 1087 -303 1126 -301
rect 1087 -305 1122 -303
rect 910 -309 940 -305
rect 952 -309 976 -305
rect 895 -315 925 -313
rect 899 -317 925 -315
rect 822 -332 826 -324
rect 822 -336 827 -332
rect 831 -336 848 -332
rect 852 -336 856 -332
rect 912 -344 917 -317
rect 952 -324 956 -309
rect 922 -336 926 -328
rect 920 -340 927 -336
rect 931 -340 948 -336
rect 952 -340 957 -336
rect 912 -348 967 -344
rect 737 -353 772 -349
rect 784 -353 804 -349
rect 727 -361 757 -357
rect 784 -368 788 -353
rect 962 -357 967 -348
rect 972 -349 976 -309
rect 1035 -313 1060 -309
rect 988 -318 994 -314
rect 998 -318 1013 -314
rect 1017 -318 1025 -314
rect 989 -328 993 -318
rect 1019 -328 1023 -318
rect 1004 -341 1008 -332
rect 1004 -345 1023 -341
rect 1019 -349 1023 -345
rect 1035 -349 1039 -313
rect 1087 -320 1091 -305
rect 1163 -307 1185 -305
rect 1198 -305 1203 -266
rect 1269 -270 1295 -266
rect 1307 -270 1327 -266
rect 1343 -270 1350 -266
rect 1354 -270 1369 -266
rect 1373 -270 1383 -266
rect 1206 -274 1215 -270
rect 1219 -274 1234 -270
rect 1238 -274 1243 -270
rect 1210 -284 1214 -274
rect 1240 -284 1244 -274
rect 1260 -278 1280 -274
rect 1225 -297 1229 -288
rect 1225 -301 1244 -297
rect 1240 -305 1244 -301
rect 1260 -305 1264 -278
rect 1307 -285 1311 -270
rect 1277 -297 1281 -289
rect 1275 -301 1282 -297
rect 1286 -301 1303 -297
rect 1307 -301 1311 -297
rect 1323 -301 1327 -270
rect 1345 -280 1349 -270
rect 1375 -280 1379 -270
rect 1360 -293 1364 -284
rect 1360 -297 1379 -293
rect 1375 -301 1379 -297
rect 1433 -301 1438 -266
rect 1504 -270 1530 -266
rect 1542 -270 1562 -266
rect 1578 -270 1585 -266
rect 1589 -270 1604 -266
rect 1608 -270 1618 -266
rect 1441 -274 1450 -270
rect 1454 -274 1469 -270
rect 1473 -274 1478 -270
rect 1445 -284 1449 -274
rect 1475 -284 1479 -274
rect 1495 -278 1515 -274
rect 1460 -297 1464 -288
rect 1460 -301 1479 -297
rect 1323 -305 1363 -301
rect 1375 -303 1438 -301
rect 1375 -305 1404 -303
rect 1189 -307 1228 -305
rect 1159 -309 1228 -307
rect 1240 -309 1264 -305
rect 1149 -315 1151 -313
rect 1155 -315 1213 -313
rect 1149 -317 1185 -315
rect 1189 -317 1213 -315
rect 1057 -332 1061 -324
rect 1057 -336 1062 -332
rect 1066 -336 1083 -332
rect 1087 -336 1091 -332
rect 1200 -344 1205 -317
rect 1240 -324 1244 -309
rect 1210 -336 1214 -328
rect 1208 -340 1215 -336
rect 1219 -340 1236 -336
rect 1240 -340 1245 -336
rect 1200 -348 1255 -344
rect 972 -353 1007 -349
rect 1019 -353 1039 -349
rect 962 -361 992 -357
rect 1019 -368 1023 -353
rect 1250 -357 1255 -348
rect 1260 -349 1264 -309
rect 1323 -313 1348 -309
rect 1276 -318 1282 -314
rect 1286 -318 1301 -314
rect 1305 -318 1313 -314
rect 1277 -328 1281 -318
rect 1307 -328 1311 -318
rect 1292 -341 1296 -332
rect 1292 -345 1311 -341
rect 1307 -349 1311 -345
rect 1323 -349 1327 -313
rect 1375 -320 1379 -305
rect 1408 -305 1438 -303
rect 1475 -305 1479 -301
rect 1495 -305 1499 -278
rect 1542 -285 1546 -270
rect 1512 -297 1516 -289
rect 1510 -301 1517 -297
rect 1521 -301 1538 -297
rect 1542 -301 1546 -297
rect 1558 -301 1562 -270
rect 1580 -280 1584 -270
rect 1610 -280 1614 -270
rect 1595 -293 1599 -284
rect 1595 -297 1614 -293
rect 1610 -301 1614 -297
rect 1558 -305 1598 -301
rect 1610 -303 1649 -301
rect 1610 -305 1645 -303
rect 1433 -309 1463 -305
rect 1475 -309 1499 -305
rect 1418 -315 1448 -313
rect 1422 -317 1448 -315
rect 1345 -332 1349 -324
rect 1345 -336 1350 -332
rect 1354 -336 1371 -332
rect 1375 -336 1379 -332
rect 1435 -344 1440 -317
rect 1475 -324 1479 -309
rect 1445 -336 1449 -328
rect 1443 -340 1450 -336
rect 1454 -340 1471 -336
rect 1475 -340 1480 -336
rect 1435 -348 1490 -344
rect 1260 -353 1295 -349
rect 1307 -353 1327 -349
rect 1250 -361 1280 -357
rect 1307 -368 1311 -353
rect 1485 -357 1490 -348
rect 1495 -349 1499 -309
rect 1558 -313 1583 -309
rect 1511 -318 1517 -314
rect 1521 -318 1536 -314
rect 1540 -318 1548 -314
rect 1512 -328 1516 -318
rect 1542 -328 1546 -318
rect 1527 -341 1531 -332
rect 1527 -345 1546 -341
rect 1542 -349 1546 -345
rect 1558 -349 1562 -313
rect 1610 -320 1614 -305
rect 1686 -307 1708 -305
rect 1721 -305 1726 -266
rect 1792 -270 1818 -266
rect 1830 -270 1850 -266
rect 1866 -270 1873 -266
rect 1877 -270 1892 -266
rect 1896 -270 1906 -266
rect 1729 -274 1738 -270
rect 1742 -274 1757 -270
rect 1761 -274 1766 -270
rect 1733 -284 1737 -274
rect 1763 -284 1767 -274
rect 1783 -278 1803 -274
rect 1748 -297 1752 -288
rect 1748 -301 1767 -297
rect 1763 -305 1767 -301
rect 1783 -305 1787 -278
rect 1830 -285 1834 -270
rect 1800 -297 1804 -289
rect 1798 -301 1805 -297
rect 1809 -301 1826 -297
rect 1830 -301 1834 -297
rect 1846 -301 1850 -270
rect 1868 -280 1872 -270
rect 1898 -280 1902 -270
rect 1883 -293 1887 -284
rect 1883 -297 1902 -293
rect 1898 -301 1902 -297
rect 1956 -301 1961 -266
rect 2027 -270 2053 -266
rect 2065 -270 2085 -266
rect 2101 -270 2108 -266
rect 2112 -270 2127 -266
rect 2131 -270 2141 -266
rect 1964 -274 1973 -270
rect 1977 -274 1992 -270
rect 1996 -274 2001 -270
rect 1968 -284 1972 -274
rect 1998 -284 2002 -274
rect 2018 -278 2038 -274
rect 1983 -297 1987 -288
rect 1983 -301 2002 -297
rect 1846 -305 1886 -301
rect 1898 -303 1961 -301
rect 1898 -305 1927 -303
rect 1712 -307 1751 -305
rect 1682 -309 1751 -307
rect 1763 -309 1787 -305
rect 1672 -315 1674 -313
rect 1678 -315 1736 -313
rect 1672 -317 1708 -315
rect 1712 -317 1736 -315
rect 1580 -332 1584 -324
rect 1580 -336 1585 -332
rect 1589 -336 1606 -332
rect 1610 -336 1614 -332
rect 1723 -344 1728 -317
rect 1763 -324 1767 -309
rect 1733 -336 1737 -328
rect 1731 -340 1738 -336
rect 1742 -340 1759 -336
rect 1763 -340 1768 -336
rect 1723 -348 1778 -344
rect 1495 -353 1530 -349
rect 1542 -353 1562 -349
rect 1485 -361 1515 -357
rect 1542 -368 1546 -353
rect 1773 -357 1778 -348
rect 1783 -349 1787 -309
rect 1846 -313 1871 -309
rect 1799 -318 1805 -314
rect 1809 -318 1824 -314
rect 1828 -318 1836 -314
rect 1800 -328 1804 -318
rect 1830 -328 1834 -318
rect 1815 -341 1819 -332
rect 1815 -345 1834 -341
rect 1830 -349 1834 -345
rect 1846 -349 1850 -313
rect 1898 -320 1902 -305
rect 1931 -305 1961 -303
rect 1998 -305 2002 -301
rect 2018 -305 2022 -278
rect 2065 -285 2069 -270
rect 2035 -297 2039 -289
rect 2033 -301 2040 -297
rect 2044 -301 2061 -297
rect 2065 -301 2069 -297
rect 2081 -301 2085 -270
rect 2103 -280 2107 -270
rect 2133 -280 2137 -270
rect 2118 -293 2122 -284
rect 2118 -297 2137 -293
rect 2133 -301 2137 -297
rect 2081 -305 2121 -301
rect 2133 -303 2172 -301
rect 2133 -305 2168 -303
rect 1956 -309 1986 -305
rect 1998 -309 2022 -305
rect 1941 -315 1971 -313
rect 1945 -317 1971 -315
rect 1868 -332 1872 -324
rect 1868 -336 1873 -332
rect 1877 -336 1894 -332
rect 1898 -336 1902 -332
rect 1958 -344 1963 -317
rect 1998 -324 2002 -309
rect 1968 -336 1972 -328
rect 1966 -340 1973 -336
rect 1977 -340 1994 -336
rect 1998 -340 2003 -336
rect 1958 -348 2013 -344
rect 1783 -353 1818 -349
rect 1830 -353 1850 -349
rect 1773 -361 1803 -357
rect 1830 -368 1834 -353
rect 2008 -357 2013 -348
rect 2018 -349 2022 -309
rect 2081 -313 2106 -309
rect 2034 -318 2040 -314
rect 2044 -318 2059 -314
rect 2063 -318 2071 -314
rect 2035 -328 2039 -318
rect 2065 -328 2069 -318
rect 2050 -341 2054 -332
rect 2050 -345 2069 -341
rect 2065 -349 2069 -345
rect 2081 -349 2085 -313
rect 2133 -320 2137 -305
rect 2209 -307 2231 -305
rect 2244 -305 2249 -266
rect 2315 -270 2341 -266
rect 2353 -270 2373 -266
rect 2389 -270 2396 -266
rect 2400 -270 2415 -266
rect 2419 -270 2429 -266
rect 2252 -274 2261 -270
rect 2265 -274 2280 -270
rect 2284 -274 2289 -270
rect 2256 -284 2260 -274
rect 2286 -284 2290 -274
rect 2306 -278 2326 -274
rect 2271 -297 2275 -288
rect 2271 -301 2290 -297
rect 2286 -305 2290 -301
rect 2306 -305 2310 -278
rect 2353 -285 2357 -270
rect 2323 -297 2327 -289
rect 2321 -301 2328 -297
rect 2332 -301 2349 -297
rect 2353 -301 2357 -297
rect 2369 -301 2373 -270
rect 2391 -280 2395 -270
rect 2421 -280 2425 -270
rect 2406 -293 2410 -284
rect 2406 -297 2425 -293
rect 2421 -301 2425 -297
rect 2479 -301 2484 -266
rect 2550 -270 2576 -266
rect 2588 -270 2608 -266
rect 2624 -270 2631 -266
rect 2635 -270 2650 -266
rect 2654 -270 2664 -266
rect 2487 -274 2496 -270
rect 2500 -274 2515 -270
rect 2519 -274 2524 -270
rect 2491 -284 2495 -274
rect 2521 -284 2525 -274
rect 2541 -278 2561 -274
rect 2506 -297 2510 -288
rect 2506 -301 2525 -297
rect 2369 -305 2409 -301
rect 2421 -303 2484 -301
rect 2421 -305 2450 -303
rect 2235 -307 2274 -305
rect 2205 -309 2274 -307
rect 2286 -309 2310 -305
rect 2195 -315 2197 -313
rect 2201 -315 2259 -313
rect 2195 -317 2231 -315
rect 2235 -317 2259 -315
rect 2103 -332 2107 -324
rect 2103 -336 2108 -332
rect 2112 -336 2129 -332
rect 2133 -336 2137 -332
rect 2246 -344 2251 -317
rect 2286 -324 2290 -309
rect 2256 -336 2260 -328
rect 2254 -340 2261 -336
rect 2265 -340 2282 -336
rect 2286 -340 2291 -336
rect 2246 -348 2301 -344
rect 2018 -353 2053 -349
rect 2065 -353 2085 -349
rect 2008 -361 2038 -357
rect 2065 -368 2069 -353
rect 2296 -357 2301 -348
rect 2306 -349 2310 -309
rect 2369 -313 2394 -309
rect 2322 -318 2328 -314
rect 2332 -318 2347 -314
rect 2351 -318 2359 -314
rect 2323 -328 2327 -318
rect 2353 -328 2357 -318
rect 2338 -341 2342 -332
rect 2338 -345 2357 -341
rect 2353 -349 2357 -345
rect 2369 -349 2373 -313
rect 2421 -320 2425 -305
rect 2454 -305 2484 -303
rect 2521 -305 2525 -301
rect 2541 -305 2545 -278
rect 2588 -285 2592 -270
rect 2558 -297 2562 -289
rect 2556 -301 2563 -297
rect 2567 -301 2584 -297
rect 2588 -301 2592 -297
rect 2604 -301 2608 -270
rect 2626 -280 2630 -270
rect 2656 -280 2660 -270
rect 2641 -293 2645 -284
rect 2641 -297 2660 -293
rect 2656 -301 2660 -297
rect 2604 -305 2644 -301
rect 2656 -303 2695 -301
rect 2656 -305 2691 -303
rect 2479 -309 2509 -305
rect 2521 -309 2545 -305
rect 2464 -315 2494 -313
rect 2468 -317 2494 -315
rect 2391 -332 2395 -324
rect 2391 -336 2396 -332
rect 2400 -336 2417 -332
rect 2421 -336 2425 -332
rect 2481 -344 2486 -317
rect 2521 -324 2525 -309
rect 2491 -336 2495 -328
rect 2489 -340 2496 -336
rect 2500 -340 2517 -336
rect 2521 -340 2526 -336
rect 2481 -348 2536 -344
rect 2306 -353 2341 -349
rect 2353 -353 2373 -349
rect 2296 -361 2326 -357
rect 2353 -368 2357 -353
rect 2531 -357 2536 -348
rect 2541 -349 2545 -309
rect 2604 -313 2629 -309
rect 2557 -318 2563 -314
rect 2567 -318 2582 -314
rect 2586 -318 2594 -314
rect 2558 -328 2562 -318
rect 2588 -328 2592 -318
rect 2573 -341 2577 -332
rect 2573 -345 2592 -341
rect 2588 -349 2592 -345
rect 2604 -349 2608 -313
rect 2656 -320 2660 -305
rect 2626 -332 2630 -324
rect 2626 -336 2631 -332
rect 2635 -336 2652 -332
rect 2656 -336 2660 -332
rect 2541 -353 2576 -349
rect 2588 -353 2608 -349
rect 2531 -361 2561 -357
rect 2588 -368 2592 -353
rect 721 -382 732 -380
rect 754 -380 758 -372
rect 736 -382 759 -380
rect 721 -384 759 -382
rect 763 -384 780 -380
rect 784 -382 792 -380
rect 796 -382 816 -380
rect 820 -382 967 -380
rect 989 -380 993 -372
rect 971 -382 994 -380
rect 784 -384 994 -382
rect 998 -384 1015 -380
rect 1019 -382 1027 -380
rect 1031 -382 1051 -380
rect 1055 -382 1119 -380
rect 1019 -384 1105 -382
rect 1109 -384 1119 -382
rect 1244 -382 1255 -380
rect 1277 -380 1281 -372
rect 1259 -382 1282 -380
rect 1244 -384 1282 -382
rect 1286 -384 1303 -380
rect 1307 -382 1315 -380
rect 1319 -382 1339 -380
rect 1343 -382 1490 -380
rect 1512 -380 1516 -372
rect 1494 -382 1517 -380
rect 1307 -384 1517 -382
rect 1521 -384 1538 -380
rect 1542 -382 1550 -380
rect 1554 -382 1574 -380
rect 1578 -382 1642 -380
rect 1542 -384 1628 -382
rect 1632 -384 1642 -382
rect 1767 -382 1778 -380
rect 1800 -380 1804 -372
rect 1782 -382 1805 -380
rect 1767 -384 1805 -382
rect 1809 -384 1826 -380
rect 1830 -382 1838 -380
rect 1842 -382 1862 -380
rect 1866 -382 2013 -380
rect 2035 -380 2039 -372
rect 2017 -382 2040 -380
rect 1830 -384 2040 -382
rect 2044 -384 2061 -380
rect 2065 -382 2073 -380
rect 2077 -382 2097 -380
rect 2101 -382 2165 -380
rect 2065 -384 2151 -382
rect 2155 -384 2165 -382
rect 2290 -382 2301 -380
rect 2323 -380 2327 -372
rect 2305 -382 2328 -380
rect 2290 -384 2328 -382
rect 2332 -384 2349 -380
rect 2353 -382 2361 -380
rect 2365 -382 2385 -380
rect 2389 -382 2536 -380
rect 2558 -380 2562 -372
rect 2540 -382 2563 -380
rect 2353 -384 2563 -382
rect 2567 -384 2584 -380
rect 2588 -382 2596 -380
rect 2600 -382 2620 -380
rect 2624 -382 2688 -380
rect 2588 -384 2674 -382
rect 2678 -384 2688 -382
rect 462 -394 895 -392
rect 462 -396 869 -394
rect 873 -396 899 -394
rect 1148 -394 1418 -392
rect 1148 -396 1392 -394
rect 665 -408 673 -404
rect 677 -408 692 -404
rect 696 -408 710 -404
rect 714 -408 724 -404
rect 728 -408 925 -404
rect 929 -408 944 -404
rect 948 -408 962 -404
rect 966 -408 976 -404
rect 980 -408 1042 -404
rect 1046 -408 1061 -404
rect 1065 -408 1079 -404
rect 1083 -408 1093 -404
rect 1097 -406 1113 -404
rect 1117 -406 1119 -404
rect 1097 -408 1119 -406
rect 668 -418 672 -408
rect 698 -418 702 -408
rect 710 -418 714 -408
rect 920 -418 924 -408
rect 950 -418 954 -408
rect 962 -418 966 -408
rect 1037 -418 1041 -408
rect 1079 -418 1083 -408
rect 683 -431 687 -422
rect 683 -435 702 -431
rect 698 -439 702 -435
rect 724 -437 728 -422
rect 935 -431 939 -422
rect 976 -431 980 -422
rect 887 -435 927 -431
rect 935 -435 954 -431
rect 698 -443 714 -439
rect 724 -441 730 -437
rect 923 -439 927 -435
rect 950 -439 954 -435
rect 976 -435 1056 -431
rect 698 -458 702 -443
rect 724 -458 728 -441
rect 923 -443 938 -439
rect 950 -443 966 -439
rect 875 -451 923 -447
rect 950 -458 954 -443
rect 976 -458 980 -435
rect 1067 -439 1071 -422
rect 1093 -437 1097 -422
rect 1148 -437 1152 -396
rect 1396 -396 1422 -394
rect 1671 -394 1941 -392
rect 1671 -396 1915 -394
rect 1188 -408 1196 -404
rect 1200 -408 1215 -404
rect 1219 -408 1233 -404
rect 1237 -408 1247 -404
rect 1251 -408 1448 -404
rect 1452 -408 1467 -404
rect 1471 -408 1485 -404
rect 1489 -408 1499 -404
rect 1503 -408 1565 -404
rect 1569 -408 1584 -404
rect 1588 -408 1602 -404
rect 1606 -408 1616 -404
rect 1620 -406 1636 -404
rect 1640 -406 1642 -404
rect 1620 -408 1642 -406
rect 1191 -418 1195 -408
rect 1221 -418 1225 -408
rect 1233 -418 1237 -408
rect 1443 -418 1447 -408
rect 1473 -418 1477 -408
rect 1485 -418 1489 -408
rect 1560 -418 1564 -408
rect 1602 -418 1606 -408
rect 1206 -431 1210 -422
rect 1206 -435 1225 -431
rect 1051 -443 1083 -439
rect 1093 -441 1152 -437
rect 1221 -439 1225 -435
rect 1247 -437 1251 -422
rect 1458 -431 1462 -422
rect 1499 -431 1503 -422
rect 1410 -435 1450 -431
rect 1458 -435 1477 -431
rect 1033 -451 1040 -447
rect 1051 -458 1055 -443
rect 1093 -458 1097 -441
rect 1221 -443 1237 -439
rect 1247 -441 1253 -437
rect 1446 -439 1450 -435
rect 1473 -439 1477 -435
rect 1499 -435 1579 -431
rect 1221 -458 1225 -443
rect 1247 -458 1251 -441
rect 1446 -443 1461 -439
rect 1473 -443 1489 -439
rect 1398 -451 1446 -447
rect 1473 -458 1477 -443
rect 1499 -458 1503 -435
rect 1590 -439 1594 -422
rect 1616 -437 1620 -422
rect 1671 -437 1675 -396
rect 1919 -396 1945 -394
rect 2194 -394 2464 -392
rect 2194 -396 2438 -394
rect 1711 -408 1719 -404
rect 1723 -408 1738 -404
rect 1742 -408 1756 -404
rect 1760 -408 1770 -404
rect 1774 -408 1971 -404
rect 1975 -408 1990 -404
rect 1994 -408 2008 -404
rect 2012 -408 2022 -404
rect 2026 -408 2088 -404
rect 2092 -408 2107 -404
rect 2111 -408 2125 -404
rect 2129 -408 2139 -404
rect 2143 -406 2159 -404
rect 2163 -406 2165 -404
rect 2143 -408 2165 -406
rect 1714 -418 1718 -408
rect 1744 -418 1748 -408
rect 1756 -418 1760 -408
rect 1966 -418 1970 -408
rect 1996 -418 2000 -408
rect 2008 -418 2012 -408
rect 2083 -418 2087 -408
rect 2125 -418 2129 -408
rect 1729 -431 1733 -422
rect 1729 -435 1748 -431
rect 1574 -443 1606 -439
rect 1616 -441 1675 -437
rect 1744 -439 1748 -435
rect 1770 -437 1774 -422
rect 1981 -431 1985 -422
rect 2022 -431 2026 -422
rect 1933 -435 1973 -431
rect 1981 -435 2000 -431
rect 1556 -451 1563 -447
rect 1574 -458 1578 -443
rect 1616 -458 1620 -441
rect 1744 -443 1760 -439
rect 1770 -441 1776 -437
rect 1969 -439 1973 -435
rect 1996 -439 2000 -435
rect 2022 -435 2102 -431
rect 1744 -458 1748 -443
rect 1770 -458 1774 -441
rect 1969 -443 1984 -439
rect 1996 -443 2012 -439
rect 1921 -451 1969 -447
rect 1996 -458 2000 -443
rect 2022 -458 2026 -435
rect 2113 -439 2117 -422
rect 2139 -437 2143 -422
rect 2194 -437 2198 -396
rect 2442 -396 2468 -394
rect 2234 -408 2242 -404
rect 2246 -408 2261 -404
rect 2265 -408 2279 -404
rect 2283 -408 2293 -404
rect 2297 -408 2494 -404
rect 2498 -408 2513 -404
rect 2517 -408 2531 -404
rect 2535 -408 2545 -404
rect 2549 -408 2611 -404
rect 2615 -408 2630 -404
rect 2634 -408 2648 -404
rect 2652 -408 2662 -404
rect 2666 -406 2682 -404
rect 2686 -406 2688 -404
rect 2666 -408 2688 -406
rect 2237 -418 2241 -408
rect 2267 -418 2271 -408
rect 2279 -418 2283 -408
rect 2489 -418 2493 -408
rect 2519 -418 2523 -408
rect 2531 -418 2535 -408
rect 2606 -418 2610 -408
rect 2648 -418 2652 -408
rect 2252 -431 2256 -422
rect 2252 -435 2271 -431
rect 2097 -443 2129 -439
rect 2139 -441 2198 -437
rect 2267 -439 2271 -435
rect 2293 -437 2297 -422
rect 2504 -431 2508 -422
rect 2545 -431 2549 -422
rect 2456 -435 2496 -431
rect 2504 -435 2523 -431
rect 2079 -451 2086 -447
rect 2097 -458 2101 -443
rect 2139 -458 2143 -441
rect 2267 -443 2283 -439
rect 2293 -441 2299 -437
rect 2492 -439 2496 -435
rect 2519 -439 2523 -435
rect 2545 -435 2625 -431
rect 2267 -458 2271 -443
rect 2293 -458 2297 -441
rect 2492 -443 2507 -439
rect 2519 -443 2535 -439
rect 2444 -451 2492 -447
rect 2519 -458 2523 -443
rect 2545 -458 2549 -435
rect 2636 -439 2640 -422
rect 2662 -437 2666 -422
rect 2620 -443 2652 -439
rect 2662 -441 2706 -437
rect 2602 -451 2609 -447
rect 2620 -458 2624 -443
rect 2662 -458 2666 -441
rect 668 -470 672 -462
rect 710 -470 714 -462
rect 920 -470 924 -462
rect 962 -470 966 -462
rect 1037 -470 1041 -462
rect 1067 -470 1071 -462
rect 1079 -470 1083 -462
rect 618 -472 673 -470
rect 614 -474 673 -472
rect 677 -474 694 -470
rect 698 -474 710 -470
rect 714 -474 725 -470
rect 729 -474 925 -470
rect 929 -474 946 -470
rect 950 -474 962 -470
rect 966 -474 977 -470
rect 981 -474 1042 -470
rect 1046 -474 1063 -470
rect 1067 -474 1079 -470
rect 1083 -474 1094 -470
rect 1098 -472 1105 -470
rect 1191 -470 1195 -462
rect 1233 -470 1237 -462
rect 1443 -470 1447 -462
rect 1485 -470 1489 -462
rect 1560 -470 1564 -462
rect 1590 -470 1594 -462
rect 1602 -470 1606 -462
rect 1109 -472 1196 -470
rect 1098 -474 1196 -472
rect 1200 -474 1217 -470
rect 1221 -474 1233 -470
rect 1237 -474 1248 -470
rect 1252 -474 1448 -470
rect 1452 -474 1469 -470
rect 1473 -474 1485 -470
rect 1489 -474 1500 -470
rect 1504 -474 1565 -470
rect 1569 -474 1586 -470
rect 1590 -474 1602 -470
rect 1606 -474 1617 -470
rect 1621 -472 1628 -470
rect 1714 -470 1718 -462
rect 1756 -470 1760 -462
rect 1966 -470 1970 -462
rect 2008 -470 2012 -462
rect 2083 -470 2087 -462
rect 2113 -470 2117 -462
rect 2125 -470 2129 -462
rect 1632 -472 1719 -470
rect 1621 -474 1719 -472
rect 1723 -474 1740 -470
rect 1744 -474 1756 -470
rect 1760 -474 1771 -470
rect 1775 -474 1971 -470
rect 1975 -474 1992 -470
rect 1996 -474 2008 -470
rect 2012 -474 2023 -470
rect 2027 -474 2088 -470
rect 2092 -474 2109 -470
rect 2113 -474 2125 -470
rect 2129 -474 2140 -470
rect 2144 -472 2151 -470
rect 2237 -470 2241 -462
rect 2279 -470 2283 -462
rect 2489 -470 2493 -462
rect 2531 -470 2535 -462
rect 2606 -470 2610 -462
rect 2636 -470 2640 -462
rect 2648 -470 2652 -462
rect 2155 -472 2242 -470
rect 2144 -474 2242 -472
rect 2246 -474 2263 -470
rect 2267 -474 2279 -470
rect 2283 -474 2294 -470
rect 2298 -474 2494 -470
rect 2498 -474 2515 -470
rect 2519 -474 2531 -470
rect 2535 -474 2546 -470
rect 2550 -474 2611 -470
rect 2615 -474 2632 -470
rect 2636 -474 2648 -470
rect 2652 -474 2663 -470
rect 2667 -472 2674 -470
rect 2678 -472 2706 -470
rect 2667 -474 2706 -472
<< metal2 >>
rect 135 1536 192 1540
rect 188 1339 192 1536
rect 756 1351 891 1355
rect 1068 1351 1172 1355
rect 90 1335 192 1339
rect 409 1338 548 1341
rect 90 1190 94 1335
rect 397 1337 548 1338
rect 756 1340 760 1351
rect 397 1334 413 1337
rect 743 1336 760 1340
rect 1038 1312 1055 1316
rect 1168 1311 1172 1351
rect 1168 1307 1300 1311
rect 367 1295 384 1299
rect 713 1297 730 1301
rect 761 1285 894 1289
rect 1069 1285 1080 1289
rect 761 1274 765 1285
rect 411 1272 547 1274
rect 400 1270 547 1272
rect 744 1270 765 1274
rect 400 1268 415 1270
rect 1076 1245 1080 1285
rect 1368 1268 1385 1272
rect 1076 1241 1300 1245
rect 1065 1206 1332 1209
rect 958 1205 986 1206
rect 712 1202 986 1205
rect 1028 1205 1332 1206
rect 1374 1205 1392 1209
rect 1028 1202 1069 1205
rect 712 1201 962 1202
rect 600 1199 628 1201
rect 360 1197 628 1199
rect 670 1200 688 1201
rect 712 1200 716 1201
rect 670 1197 716 1200
rect 360 1195 604 1197
rect 256 1190 284 1193
rect 90 1189 284 1190
rect 326 1190 344 1193
rect 360 1190 364 1195
rect 326 1189 364 1190
rect 90 1186 260 1189
rect 90 1041 94 1186
rect 256 1145 260 1186
rect 340 1186 364 1189
rect 340 1149 344 1186
rect 600 1153 604 1195
rect 684 1196 716 1197
rect 684 1157 688 1196
rect 958 1158 962 1201
rect 1042 1162 1046 1202
rect 1042 1158 1052 1162
rect 1304 1161 1308 1205
rect 1388 1165 1392 1205
rect 1388 1161 1398 1165
rect 684 1153 694 1157
rect 910 1154 918 1158
rect 960 1154 962 1158
rect 1256 1157 1264 1161
rect 1306 1157 1308 1161
rect 552 1149 560 1153
rect 602 1149 604 1153
rect 340 1145 350 1149
rect 208 1141 216 1145
rect 258 1141 260 1145
rect 208 1071 212 1141
rect 263 1123 282 1127
rect 327 1123 346 1127
rect 263 1079 267 1123
rect 260 1075 267 1079
rect 279 1106 284 1110
rect 279 1071 283 1106
rect 342 1083 346 1123
rect 342 1079 352 1083
rect 552 1079 556 1149
rect 607 1131 626 1135
rect 671 1131 690 1135
rect 607 1087 611 1131
rect 604 1083 611 1087
rect 623 1114 628 1118
rect 623 1079 627 1114
rect 686 1091 690 1131
rect 686 1087 696 1091
rect 208 1067 283 1071
rect 350 1052 354 1079
rect 552 1075 627 1079
rect 694 1057 698 1087
rect 910 1084 914 1154
rect 965 1136 984 1140
rect 1029 1136 1048 1140
rect 965 1092 969 1136
rect 962 1088 969 1092
rect 981 1119 986 1123
rect 981 1084 985 1119
rect 1044 1096 1048 1136
rect 1044 1092 1054 1096
rect 910 1080 985 1084
rect 1052 1060 1056 1092
rect 1256 1087 1260 1157
rect 1311 1139 1330 1143
rect 1375 1139 1394 1143
rect 1311 1095 1315 1139
rect 1308 1091 1315 1095
rect 1327 1122 1332 1126
rect 1327 1087 1331 1122
rect 1390 1099 1394 1139
rect 1390 1095 1400 1099
rect 1256 1083 1331 1087
rect 1398 1060 1402 1095
rect 1052 1057 1330 1060
rect 694 1053 984 1057
rect 1030 1056 1330 1057
rect 1376 1056 1402 1060
rect 1030 1053 1056 1056
rect 694 1052 698 1053
rect 350 1048 626 1052
rect 672 1048 698 1052
rect 350 1044 354 1048
rect -130 1037 -101 1041
rect 1 1037 117 1041
rect 328 1040 354 1044
rect -130 877 -126 1037
rect 1 970 97 974
rect 93 901 97 970
rect 113 968 117 1037
rect 1197 1027 1308 1031
rect 1197 988 1201 1027
rect 1376 988 1393 992
rect 726 984 881 988
rect 1060 984 1201 988
rect 395 972 521 976
rect 726 975 730 984
rect 113 964 178 968
rect 395 967 399 972
rect 715 971 730 975
rect 383 963 399 967
rect 1189 961 1308 965
rect 1030 945 1047 949
rect 685 932 702 936
rect 353 924 370 928
rect 1189 922 1193 961
rect 746 918 885 922
rect 1061 918 1193 922
rect 746 909 750 918
rect 393 905 521 909
rect 716 905 750 909
rect 393 901 397 905
rect 93 897 178 901
rect 383 897 397 901
rect -130 873 -49 877
rect -97 152 -93 873
rect 93 810 97 897
rect 82 806 97 810
rect -45 274 -41 287
rect 27 274 31 775
rect -45 270 31 274
rect 111 279 115 287
rect 111 275 129 279
rect -45 203 -41 270
rect -47 199 -41 203
rect -806 148 -800 152
rect -168 148 -93 152
rect -806 -27 -802 148
rect -97 103 -93 148
rect -82 133 -76 137
rect -82 103 -78 133
rect -45 119 -41 199
rect -47 115 -41 119
rect 111 203 115 275
rect 201 209 220 213
rect 111 199 131 203
rect 111 127 115 199
rect 216 137 220 209
rect 203 133 230 137
rect 111 123 133 127
rect -97 99 -78 103
rect -82 53 -78 99
rect -82 49 -76 53
rect 111 51 115 123
rect 216 61 220 133
rect 205 57 220 61
rect -82 -24 -78 49
rect 111 47 135 51
rect 216 -15 220 57
rect 207 -19 220 -15
rect -806 -31 -622 -27
rect 216 -24 220 -19
rect 262 19 264 23
rect 262 -26 266 19
rect 229 -30 266 -26
rect 262 -460 266 -30
rect 455 -86 459 -53
rect 968 -86 972 -53
rect 1474 -86 1478 -53
rect 1998 -86 2002 -53
rect 457 -90 467 -86
rect 970 -90 980 -86
rect 1476 -90 1486 -86
rect 2000 -90 2010 -86
rect 463 -130 467 -90
rect 463 -134 482 -130
rect 459 -156 469 -152
rect 465 -194 469 -156
rect 525 -194 529 -113
rect 976 -130 980 -90
rect 976 -134 995 -130
rect 549 -152 551 -148
rect 549 -194 553 -152
rect 972 -156 982 -152
rect 978 -194 982 -156
rect 1038 -194 1042 -113
rect 1482 -130 1486 -90
rect 1482 -134 1501 -130
rect 1062 -152 1064 -148
rect 1062 -194 1066 -152
rect 1478 -156 1488 -152
rect 1484 -194 1488 -156
rect 1544 -194 1548 -113
rect 2006 -130 2010 -90
rect 2006 -134 2025 -130
rect 1568 -152 1570 -148
rect 1568 -194 1572 -152
rect 2002 -156 2012 -152
rect 2008 -194 2012 -156
rect 2068 -194 2072 -113
rect 2092 -152 2094 -148
rect 2092 -194 2096 -152
rect 590 -340 594 -202
rect 722 -270 726 -237
rect 957 -270 961 -237
rect 724 -274 734 -270
rect 959 -274 969 -270
rect 730 -314 734 -274
rect 730 -318 749 -314
rect 726 -340 736 -336
rect 590 -344 618 -340
rect 614 -460 618 -344
rect 732 -378 736 -340
rect 792 -378 796 -297
rect 965 -314 969 -274
rect 965 -318 984 -314
rect 816 -336 818 -332
rect 816 -378 820 -336
rect 961 -340 971 -336
rect 967 -378 971 -340
rect 1027 -378 1031 -297
rect 1051 -336 1053 -332
rect 1051 -378 1055 -336
rect 262 -464 618 -460
rect 614 -468 618 -464
rect 1105 -468 1109 -386
rect 1113 -402 1117 -237
rect 1245 -270 1249 -237
rect 1480 -270 1484 -237
rect 1247 -274 1257 -270
rect 1482 -274 1492 -270
rect 1253 -314 1257 -274
rect 1253 -318 1272 -314
rect 1249 -340 1259 -336
rect 1255 -378 1259 -340
rect 1315 -378 1319 -297
rect 1488 -314 1492 -274
rect 1488 -318 1507 -314
rect 1339 -336 1341 -332
rect 1339 -378 1343 -336
rect 1484 -340 1494 -336
rect 1490 -378 1494 -340
rect 1550 -378 1554 -297
rect 1574 -336 1576 -332
rect 1574 -378 1578 -336
rect 1628 -468 1632 -386
rect 1636 -402 1640 -237
rect 1768 -270 1772 -237
rect 2003 -270 2007 -237
rect 1770 -274 1780 -270
rect 2005 -274 2015 -270
rect 1776 -314 1780 -274
rect 1776 -318 1795 -314
rect 1772 -340 1782 -336
rect 1778 -378 1782 -340
rect 1838 -378 1842 -297
rect 2011 -314 2015 -274
rect 2011 -318 2030 -314
rect 1862 -336 1864 -332
rect 1862 -378 1866 -336
rect 2007 -340 2017 -336
rect 2013 -378 2017 -340
rect 2073 -378 2077 -297
rect 2097 -336 2099 -332
rect 2097 -378 2101 -336
rect 2151 -468 2155 -386
rect 2159 -402 2163 -237
rect 2291 -270 2295 -237
rect 2526 -270 2530 -237
rect 2293 -274 2303 -270
rect 2528 -274 2538 -270
rect 2299 -314 2303 -274
rect 2299 -318 2318 -314
rect 2295 -340 2305 -336
rect 2301 -378 2305 -340
rect 2361 -378 2365 -297
rect 2534 -314 2538 -274
rect 2534 -318 2553 -314
rect 2385 -336 2387 -332
rect 2385 -378 2389 -336
rect 2530 -340 2540 -336
rect 2536 -378 2540 -340
rect 2596 -378 2600 -297
rect 2620 -336 2622 -332
rect 2620 -378 2624 -336
rect 2674 -468 2678 -386
rect 2682 -402 2686 -237
<< ntransistor >>
rect 18 1522 20 1530
rect 44 1522 47 1530
rect 68 1522 71 1530
rect 94 1522 97 1530
rect 118 1522 121 1530
rect 907 1337 909 1345
rect 933 1337 936 1345
rect 948 1337 951 1345
rect 206 1321 208 1329
rect 232 1321 235 1329
rect 247 1321 250 1329
rect 262 1321 265 1329
rect 277 1321 280 1329
rect 313 1320 315 1328
rect 339 1320 342 1328
rect 354 1320 357 1328
rect 381 1320 383 1328
rect 563 1323 565 1331
rect 589 1323 592 1331
rect 604 1323 607 1331
rect 619 1323 622 1331
rect 659 1322 661 1330
rect 685 1322 688 1330
rect 700 1322 703 1330
rect 727 1322 729 1330
rect 984 1337 986 1345
rect 1010 1337 1013 1345
rect 1025 1337 1028 1345
rect 1052 1337 1054 1345
rect 1314 1293 1316 1301
rect 1340 1293 1343 1301
rect 1355 1293 1358 1301
rect 1382 1293 1384 1301
rect 640 1183 643 1191
rect 655 1183 658 1191
rect 998 1188 1001 1196
rect 1013 1188 1016 1196
rect 1344 1191 1347 1199
rect 1359 1191 1362 1199
rect 296 1175 299 1183
rect 311 1175 314 1183
rect 228 1127 231 1135
rect 243 1127 246 1135
rect 363 1131 366 1139
rect 378 1131 381 1139
rect 572 1135 575 1143
rect 587 1135 590 1143
rect 707 1139 710 1147
rect 722 1139 725 1147
rect 930 1140 933 1148
rect 945 1140 948 1148
rect 1065 1144 1068 1152
rect 1080 1144 1083 1152
rect 171 1118 173 1126
rect -87 1023 -85 1031
rect -61 1023 -58 1031
rect -46 1023 -43 1031
rect -31 1023 -28 1031
rect -16 1023 -13 1031
rect 515 1126 517 1134
rect 296 1092 299 1100
rect 311 1092 314 1100
rect 873 1131 875 1139
rect 640 1100 643 1108
rect 655 1100 658 1108
rect 1276 1143 1279 1151
rect 1291 1143 1294 1151
rect 1411 1147 1414 1155
rect 1426 1147 1429 1155
rect 998 1105 1001 1113
rect 1013 1105 1016 1113
rect 1219 1134 1221 1142
rect 1344 1108 1347 1116
rect 1359 1108 1362 1116
rect 1322 1013 1324 1021
rect 1348 1013 1351 1021
rect 1363 1013 1366 1021
rect 1390 1013 1392 1021
rect 899 970 901 978
rect 925 970 928 978
rect 940 970 943 978
rect 192 950 194 958
rect 218 950 221 958
rect 233 950 236 958
rect 248 950 251 958
rect 263 950 266 958
rect 535 958 537 966
rect 561 958 564 966
rect 576 958 579 966
rect 591 958 594 966
rect 299 949 301 957
rect 325 949 328 957
rect 340 949 343 957
rect 367 949 369 957
rect 631 957 633 965
rect 657 957 660 965
rect 672 957 675 965
rect 699 957 701 965
rect 976 970 978 978
rect 1002 970 1005 978
rect 1017 970 1020 978
rect 1044 970 1046 978
rect -35 859 -33 867
rect -9 859 -6 867
rect 15 859 18 867
rect 41 859 44 867
rect 65 859 68 867
rect -784 158 -781 166
rect -769 158 -766 166
rect -742 158 -740 166
rect -707 158 -704 166
rect -692 158 -689 166
rect -665 158 -663 166
rect -630 158 -627 166
rect -615 158 -612 166
rect -588 158 -586 166
rect -553 158 -550 166
rect -538 158 -535 166
rect -511 158 -509 166
rect -476 158 -473 166
rect -461 158 -458 166
rect -434 158 -432 166
rect -399 158 -396 166
rect -384 158 -381 166
rect -357 158 -355 166
rect -322 158 -319 166
rect -307 158 -304 166
rect -280 158 -278 166
rect -245 158 -242 166
rect -230 158 -227 166
rect -203 158 -201 166
rect -63 143 -61 151
rect -63 59 -61 67
rect 143 219 146 227
rect 158 219 161 227
rect 185 219 187 227
rect 145 143 148 151
rect 160 143 163 151
rect 187 143 189 151
rect 291 143 294 151
rect 306 143 309 151
rect 333 143 335 151
rect 461 143 464 151
rect 476 143 479 151
rect 503 143 505 151
rect 849 143 852 151
rect 864 143 867 151
rect 891 143 893 151
rect 1019 143 1022 151
rect 1034 143 1037 151
rect 1061 143 1063 151
rect 1354 143 1357 151
rect 1369 143 1372 151
rect 1396 143 1398 151
rect 1524 143 1527 151
rect 1539 143 1542 151
rect 1566 143 1568 151
rect 1878 143 1881 151
rect 1893 143 1896 151
rect 1920 143 1922 151
rect 2048 143 2051 151
rect 2063 143 2066 151
rect 2090 143 2092 151
rect -609 -21 -606 -13
rect -594 -21 -591 -13
rect -567 -21 -565 -13
rect -532 -21 -529 -13
rect -517 -21 -514 -13
rect -490 -21 -488 -13
rect -455 -21 -452 -13
rect -440 -21 -437 -13
rect -413 -21 -411 -13
rect -378 -21 -375 -13
rect -363 -21 -360 -13
rect -336 -21 -334 -13
rect 147 67 150 75
rect 162 67 165 75
rect 189 67 191 75
rect 276 29 279 37
rect 291 29 294 37
rect 318 29 320 37
rect 398 29 401 37
rect 413 29 416 37
rect 440 29 442 37
rect 568 29 571 37
rect 583 29 586 37
rect 610 29 612 37
rect 149 -9 152 -1
rect 164 -9 167 -1
rect 191 -9 193 -1
rect 495 -107 498 -99
rect 510 -107 513 -99
rect 428 -146 431 -138
rect 443 -146 446 -138
rect 563 -142 566 -134
rect 578 -142 581 -134
rect 495 -190 498 -182
rect 510 -190 513 -182
rect 956 29 959 37
rect 971 29 974 37
rect 998 29 1000 37
rect 1126 29 1129 37
rect 1141 29 1144 37
rect 1168 29 1170 37
rect 1461 29 1464 37
rect 1476 29 1479 37
rect 1503 29 1505 37
rect 1631 29 1634 37
rect 1646 29 1649 37
rect 1673 29 1675 37
rect 1008 -107 1011 -99
rect 1023 -107 1026 -99
rect 941 -146 944 -138
rect 956 -146 959 -138
rect 1076 -142 1079 -134
rect 1091 -142 1094 -134
rect 1008 -190 1011 -182
rect 1023 -190 1026 -182
rect 762 -291 765 -283
rect 777 -291 780 -283
rect 695 -330 698 -322
rect 710 -330 713 -322
rect 830 -326 833 -318
rect 845 -326 848 -318
rect 762 -374 765 -366
rect 777 -374 780 -366
rect 676 -464 679 -456
rect 691 -464 694 -456
rect 718 -464 720 -456
rect 997 -291 1000 -283
rect 1012 -291 1015 -283
rect 930 -330 933 -322
rect 945 -330 948 -322
rect 1065 -326 1068 -318
rect 1080 -326 1083 -318
rect 997 -374 1000 -366
rect 1012 -374 1015 -366
rect 928 -464 931 -456
rect 943 -464 946 -456
rect 970 -464 972 -456
rect 1045 -464 1048 -456
rect 1060 -464 1063 -456
rect 1087 -464 1089 -456
rect 1985 29 1988 37
rect 2000 29 2003 37
rect 2027 29 2029 37
rect 2155 29 2158 37
rect 2170 29 2173 37
rect 2197 29 2199 37
rect 1514 -107 1517 -99
rect 1529 -107 1532 -99
rect 1447 -146 1450 -138
rect 1462 -146 1465 -138
rect 1582 -142 1585 -134
rect 1597 -142 1600 -134
rect 1514 -190 1517 -182
rect 1529 -190 1532 -182
rect 1285 -291 1288 -283
rect 1300 -291 1303 -283
rect 1218 -330 1221 -322
rect 1233 -330 1236 -322
rect 1353 -326 1356 -318
rect 1368 -326 1371 -318
rect 1285 -374 1288 -366
rect 1300 -374 1303 -366
rect 1199 -464 1202 -456
rect 1214 -464 1217 -456
rect 1241 -464 1243 -456
rect 1520 -291 1523 -283
rect 1535 -291 1538 -283
rect 1453 -330 1456 -322
rect 1468 -330 1471 -322
rect 1588 -326 1591 -318
rect 1603 -326 1606 -318
rect 1520 -374 1523 -366
rect 1535 -374 1538 -366
rect 1451 -464 1454 -456
rect 1466 -464 1469 -456
rect 1493 -464 1495 -456
rect 1568 -464 1571 -456
rect 1583 -464 1586 -456
rect 1610 -464 1612 -456
rect 2038 -107 2041 -99
rect 2053 -107 2056 -99
rect 1971 -146 1974 -138
rect 1986 -146 1989 -138
rect 2106 -142 2109 -134
rect 2121 -142 2124 -134
rect 2038 -190 2041 -182
rect 2053 -190 2056 -182
rect 1808 -291 1811 -283
rect 1823 -291 1826 -283
rect 1741 -330 1744 -322
rect 1756 -330 1759 -322
rect 1876 -326 1879 -318
rect 1891 -326 1894 -318
rect 1808 -374 1811 -366
rect 1823 -374 1826 -366
rect 1722 -464 1725 -456
rect 1737 -464 1740 -456
rect 1764 -464 1766 -456
rect 2043 -291 2046 -283
rect 2058 -291 2061 -283
rect 1976 -330 1979 -322
rect 1991 -330 1994 -322
rect 2111 -326 2114 -318
rect 2126 -326 2129 -318
rect 2043 -374 2046 -366
rect 2058 -374 2061 -366
rect 1974 -464 1977 -456
rect 1989 -464 1992 -456
rect 2016 -464 2018 -456
rect 2091 -464 2094 -456
rect 2106 -464 2109 -456
rect 2133 -464 2135 -456
rect 2331 -291 2334 -283
rect 2346 -291 2349 -283
rect 2264 -330 2267 -322
rect 2279 -330 2282 -322
rect 2399 -326 2402 -318
rect 2414 -326 2417 -318
rect 2331 -374 2334 -366
rect 2346 -374 2349 -366
rect 2245 -464 2248 -456
rect 2260 -464 2263 -456
rect 2287 -464 2289 -456
rect 2566 -291 2569 -283
rect 2581 -291 2584 -283
rect 2499 -330 2502 -322
rect 2514 -330 2517 -322
rect 2634 -326 2637 -318
rect 2649 -326 2652 -318
rect 2566 -374 2569 -366
rect 2581 -374 2584 -366
rect 2497 -464 2500 -456
rect 2512 -464 2515 -456
rect 2539 -464 2541 -456
rect 2614 -464 2617 -456
rect 2629 -464 2632 -456
rect 2656 -464 2658 -456
<< ptransistor >>
rect 18 1481 20 1489
rect 44 1481 47 1489
rect 68 1481 71 1489
rect 94 1481 97 1489
rect 118 1481 121 1489
rect 907 1297 909 1305
rect 933 1297 936 1305
rect 948 1297 951 1305
rect 984 1297 986 1305
rect 1010 1297 1013 1305
rect 1025 1297 1028 1305
rect 1052 1297 1054 1305
rect 206 1280 208 1288
rect 232 1280 235 1288
rect 247 1280 250 1288
rect 262 1280 265 1288
rect 277 1280 280 1288
rect 313 1280 315 1288
rect 339 1280 342 1288
rect 354 1280 357 1288
rect 381 1280 383 1288
rect 563 1282 565 1290
rect 589 1282 592 1290
rect 604 1282 607 1290
rect 619 1282 622 1290
rect 659 1282 661 1290
rect 685 1282 688 1290
rect 700 1282 703 1290
rect 727 1282 729 1290
rect 1314 1253 1316 1261
rect 1340 1253 1343 1261
rect 1355 1253 1358 1261
rect 1382 1253 1384 1261
rect 296 1135 299 1143
rect 311 1135 314 1143
rect 640 1143 643 1151
rect 655 1143 658 1151
rect 998 1148 1001 1156
rect 1013 1148 1016 1156
rect 1344 1151 1347 1159
rect 1359 1151 1362 1159
rect 171 1096 173 1104
rect 228 1087 231 1095
rect 243 1087 246 1095
rect 515 1104 517 1112
rect 363 1091 366 1099
rect 378 1091 381 1099
rect 572 1095 575 1103
rect 587 1095 590 1103
rect 873 1109 875 1117
rect 707 1099 710 1107
rect 722 1099 725 1107
rect 930 1100 933 1108
rect 945 1100 948 1108
rect 1219 1112 1221 1120
rect 1065 1104 1068 1112
rect 1080 1104 1083 1112
rect 1276 1103 1279 1111
rect 1291 1103 1294 1111
rect 1411 1107 1414 1115
rect 1426 1107 1429 1115
rect 640 1060 643 1068
rect 655 1060 658 1068
rect 998 1065 1001 1073
rect 1013 1065 1016 1073
rect 1344 1068 1347 1076
rect 1359 1068 1362 1076
rect 296 1052 299 1060
rect 311 1052 314 1060
rect -87 982 -85 990
rect -61 982 -58 990
rect -46 982 -43 990
rect -31 982 -28 990
rect -16 982 -13 990
rect 1322 973 1324 981
rect 1348 973 1351 981
rect 1363 973 1366 981
rect 1390 973 1392 981
rect 899 930 901 938
rect 925 930 928 938
rect 940 930 943 938
rect 976 930 978 938
rect 1002 930 1005 938
rect 1017 930 1020 938
rect 1044 930 1046 938
rect 535 917 537 925
rect 561 917 564 925
rect 576 917 579 925
rect 591 917 594 925
rect 631 917 633 925
rect 657 917 660 925
rect 672 917 675 925
rect 699 917 701 925
rect 192 909 194 917
rect 218 909 221 917
rect 233 909 236 917
rect 248 909 251 917
rect 263 909 266 917
rect 299 909 301 917
rect 325 909 328 917
rect 340 909 343 917
rect 367 909 369 917
rect -35 818 -33 826
rect -9 818 -6 826
rect 15 818 18 826
rect 41 818 44 826
rect 65 818 68 826
rect 143 259 146 267
rect 158 259 161 267
rect 185 259 187 267
rect -784 198 -781 206
rect -769 198 -766 206
rect -742 198 -740 206
rect -707 198 -704 206
rect -692 198 -689 206
rect -665 198 -663 206
rect -630 198 -627 206
rect -615 198 -612 206
rect -588 198 -586 206
rect -553 198 -550 206
rect -538 198 -535 206
rect -511 198 -509 206
rect -476 198 -473 206
rect -461 198 -458 206
rect -434 198 -432 206
rect -399 198 -396 206
rect -384 198 -381 206
rect -357 198 -355 206
rect -322 198 -319 206
rect -307 198 -304 206
rect -280 198 -278 206
rect -245 198 -242 206
rect -230 198 -227 206
rect -203 198 -201 206
rect -63 183 -61 191
rect -63 99 -61 107
rect 145 183 148 191
rect 160 183 163 191
rect 187 183 189 191
rect 291 183 294 191
rect 306 183 309 191
rect 333 183 335 191
rect 461 183 464 191
rect 476 183 479 191
rect 503 183 505 191
rect 849 183 852 191
rect 864 183 867 191
rect 891 183 893 191
rect 1019 183 1022 191
rect 1034 183 1037 191
rect 1061 183 1063 191
rect 1354 183 1357 191
rect 1369 183 1372 191
rect 1396 183 1398 191
rect 1524 183 1527 191
rect 1539 183 1542 191
rect 1566 183 1568 191
rect 1878 183 1881 191
rect 1893 183 1896 191
rect 1920 183 1922 191
rect 2048 183 2051 191
rect 2063 183 2066 191
rect 2090 183 2092 191
rect 147 107 150 115
rect 162 107 165 115
rect 189 107 191 115
rect -609 19 -606 27
rect -594 19 -591 27
rect -567 19 -565 27
rect -532 19 -529 27
rect -517 19 -514 27
rect -490 19 -488 27
rect -455 19 -452 27
rect -440 19 -437 27
rect -413 19 -411 27
rect -378 19 -375 27
rect -363 19 -360 27
rect -336 19 -334 27
rect 276 69 279 77
rect 291 69 294 77
rect 318 69 320 77
rect 149 31 152 39
rect 164 31 167 39
rect 191 31 193 39
rect 398 69 401 77
rect 413 69 416 77
rect 440 69 442 77
rect 568 69 571 77
rect 583 69 586 77
rect 610 69 612 77
rect 956 69 959 77
rect 971 69 974 77
rect 998 69 1000 77
rect 495 -67 498 -59
rect 510 -67 513 -59
rect 428 -106 431 -98
rect 443 -106 446 -98
rect 563 -102 566 -94
rect 578 -102 581 -94
rect 495 -150 498 -142
rect 510 -150 513 -142
rect 1126 69 1129 77
rect 1141 69 1144 77
rect 1168 69 1170 77
rect 1461 69 1464 77
rect 1476 69 1479 77
rect 1503 69 1505 77
rect 1631 69 1634 77
rect 1646 69 1649 77
rect 1673 69 1675 77
rect 1985 69 1988 77
rect 2000 69 2003 77
rect 2027 69 2029 77
rect 1008 -67 1011 -59
rect 1023 -67 1026 -59
rect 941 -106 944 -98
rect 956 -106 959 -98
rect 1076 -102 1079 -94
rect 1091 -102 1094 -94
rect 1008 -150 1011 -142
rect 1023 -150 1026 -142
rect 762 -251 765 -243
rect 777 -251 780 -243
rect 997 -251 1000 -243
rect 1012 -251 1015 -243
rect 695 -290 698 -282
rect 710 -290 713 -282
rect 830 -286 833 -278
rect 845 -286 848 -278
rect 930 -290 933 -282
rect 945 -290 948 -282
rect 762 -334 765 -326
rect 777 -334 780 -326
rect 676 -424 679 -416
rect 691 -424 694 -416
rect 718 -424 720 -416
rect 1065 -286 1068 -278
rect 1080 -286 1083 -278
rect 997 -334 1000 -326
rect 1012 -334 1015 -326
rect 928 -424 931 -416
rect 943 -424 946 -416
rect 970 -424 972 -416
rect 1045 -424 1048 -416
rect 1060 -424 1063 -416
rect 1087 -424 1089 -416
rect 2155 69 2158 77
rect 2170 69 2173 77
rect 2197 69 2199 77
rect 1514 -67 1517 -59
rect 1529 -67 1532 -59
rect 1447 -106 1450 -98
rect 1462 -106 1465 -98
rect 1582 -102 1585 -94
rect 1597 -102 1600 -94
rect 1514 -150 1517 -142
rect 1529 -150 1532 -142
rect 1285 -251 1288 -243
rect 1300 -251 1303 -243
rect 1520 -251 1523 -243
rect 1535 -251 1538 -243
rect 1218 -290 1221 -282
rect 1233 -290 1236 -282
rect 1353 -286 1356 -278
rect 1368 -286 1371 -278
rect 1453 -290 1456 -282
rect 1468 -290 1471 -282
rect 1285 -334 1288 -326
rect 1300 -334 1303 -326
rect 1199 -424 1202 -416
rect 1214 -424 1217 -416
rect 1241 -424 1243 -416
rect 1588 -286 1591 -278
rect 1603 -286 1606 -278
rect 1520 -334 1523 -326
rect 1535 -334 1538 -326
rect 1451 -424 1454 -416
rect 1466 -424 1469 -416
rect 1493 -424 1495 -416
rect 1568 -424 1571 -416
rect 1583 -424 1586 -416
rect 1610 -424 1612 -416
rect 2038 -67 2041 -59
rect 2053 -67 2056 -59
rect 1971 -106 1974 -98
rect 1986 -106 1989 -98
rect 2106 -102 2109 -94
rect 2121 -102 2124 -94
rect 2038 -150 2041 -142
rect 2053 -150 2056 -142
rect 1808 -251 1811 -243
rect 1823 -251 1826 -243
rect 2043 -251 2046 -243
rect 2058 -251 2061 -243
rect 1741 -290 1744 -282
rect 1756 -290 1759 -282
rect 1876 -286 1879 -278
rect 1891 -286 1894 -278
rect 1976 -290 1979 -282
rect 1991 -290 1994 -282
rect 1808 -334 1811 -326
rect 1823 -334 1826 -326
rect 1722 -424 1725 -416
rect 1737 -424 1740 -416
rect 1764 -424 1766 -416
rect 2111 -286 2114 -278
rect 2126 -286 2129 -278
rect 2043 -334 2046 -326
rect 2058 -334 2061 -326
rect 1974 -424 1977 -416
rect 1989 -424 1992 -416
rect 2016 -424 2018 -416
rect 2091 -424 2094 -416
rect 2106 -424 2109 -416
rect 2133 -424 2135 -416
rect 2331 -251 2334 -243
rect 2346 -251 2349 -243
rect 2566 -251 2569 -243
rect 2581 -251 2584 -243
rect 2264 -290 2267 -282
rect 2279 -290 2282 -282
rect 2399 -286 2402 -278
rect 2414 -286 2417 -278
rect 2499 -290 2502 -282
rect 2514 -290 2517 -282
rect 2331 -334 2334 -326
rect 2346 -334 2349 -326
rect 2245 -424 2248 -416
rect 2260 -424 2263 -416
rect 2287 -424 2289 -416
rect 2634 -286 2637 -278
rect 2649 -286 2652 -278
rect 2566 -334 2569 -326
rect 2581 -334 2584 -326
rect 2497 -424 2500 -416
rect 2512 -424 2515 -416
rect 2539 -424 2541 -416
rect 2614 -424 2617 -416
rect 2629 -424 2632 -416
rect 2656 -424 2658 -416
<< polycontact >>
rect 20 1504 24 1508
rect 47 1494 51 1498
rect 71 1501 75 1505
rect 97 1508 101 1512
rect 121 1515 125 1519
rect 231 1398 235 1402
rect 588 1398 592 1402
rect 1174 1400 1178 1404
rect 246 1389 250 1393
rect 831 1391 835 1395
rect 485 1381 489 1385
rect 231 1368 235 1372
rect 246 1368 250 1372
rect 588 1378 592 1382
rect 208 1304 212 1308
rect 280 1293 284 1297
rect 358 1311 362 1315
rect 315 1303 319 1307
rect 343 1303 347 1307
rect 383 1312 387 1316
rect 393 1312 397 1316
rect 446 1312 450 1316
rect 393 1295 397 1299
rect 429 1295 433 1299
rect 565 1306 569 1310
rect 592 1316 596 1320
rect 622 1295 626 1299
rect 704 1313 708 1317
rect 661 1305 665 1309
rect 689 1305 693 1309
rect 729 1314 733 1318
rect 739 1314 743 1318
rect 790 1314 794 1318
rect 909 1320 913 1324
rect 937 1320 941 1324
rect 1029 1328 1033 1332
rect 986 1320 990 1324
rect 1014 1320 1018 1324
rect 1054 1329 1058 1333
rect 1064 1329 1068 1333
rect 1148 1329 1152 1333
rect 1064 1312 1068 1316
rect 1131 1312 1135 1316
rect 739 1297 743 1301
rect 773 1297 777 1301
rect 1359 1284 1363 1288
rect 1316 1276 1320 1280
rect 1344 1276 1348 1280
rect 1384 1285 1388 1289
rect 1394 1285 1398 1289
rect 1494 1285 1498 1289
rect 1394 1268 1398 1272
rect 1477 1268 1481 1272
rect 659 1174 663 1178
rect 1017 1179 1021 1183
rect 315 1166 319 1170
rect 644 1166 648 1170
rect 300 1158 304 1162
rect 1002 1171 1006 1175
rect 1363 1182 1367 1186
rect 1348 1174 1352 1178
rect 153 1109 157 1113
rect 247 1118 251 1122
rect 382 1122 386 1126
rect 410 1122 414 1126
rect 429 1122 433 1126
rect 173 1110 177 1114
rect 232 1110 236 1114
rect 367 1114 371 1118
rect 410 1114 414 1118
rect 446 1114 450 1118
rect 591 1126 595 1130
rect 726 1130 730 1134
rect 754 1130 758 1134
rect 773 1130 777 1134
rect 517 1118 521 1122
rect 576 1118 580 1122
rect 711 1122 715 1126
rect 754 1122 758 1126
rect 790 1122 794 1126
rect 949 1131 953 1135
rect 1084 1135 1088 1139
rect 1112 1135 1116 1139
rect 1131 1135 1135 1139
rect 875 1123 879 1127
rect 934 1123 938 1127
rect 1069 1127 1073 1131
rect 1112 1127 1116 1131
rect 1148 1127 1152 1131
rect 1295 1134 1299 1138
rect 1430 1138 1434 1142
rect 1458 1138 1462 1142
rect 1477 1138 1481 1142
rect 1221 1126 1225 1130
rect 1280 1126 1284 1130
rect 659 1091 663 1095
rect 1415 1130 1419 1134
rect 1458 1130 1462 1134
rect 1494 1130 1498 1134
rect 1017 1096 1021 1100
rect 315 1083 319 1087
rect 644 1083 648 1087
rect 300 1075 304 1079
rect 1002 1088 1006 1092
rect 1363 1099 1367 1103
rect 1348 1091 1352 1095
rect -85 1006 -81 1010
rect -58 1016 -54 1020
rect -43 1009 -39 1013
rect -28 1002 -24 1006
rect -1 1016 3 1020
rect -1 1009 3 1013
rect 222 1008 226 1012
rect 485 1010 489 1014
rect -1 1002 3 1006
rect 232 999 236 1003
rect 564 999 568 1003
rect 831 1001 835 1005
rect -13 995 -9 999
rect -1 995 3 999
rect 1178 991 1182 995
rect 222 981 226 985
rect 232 981 236 985
rect 564 979 568 983
rect 194 933 198 937
rect 266 922 270 926
rect 344 940 348 944
rect 301 932 305 936
rect 329 932 333 936
rect 369 941 373 945
rect 379 941 383 945
rect 429 941 433 945
rect 379 924 383 928
rect 446 924 450 928
rect 537 941 541 945
rect 564 951 568 955
rect 594 930 598 934
rect 676 948 680 952
rect 633 940 637 944
rect 661 940 665 944
rect 701 949 705 953
rect 711 949 715 953
rect 773 949 777 953
rect 1367 1004 1371 1008
rect 1324 996 1328 1000
rect 1352 996 1356 1000
rect 1392 1005 1396 1009
rect 1402 1005 1406 1009
rect 1477 1005 1481 1009
rect 1402 988 1406 992
rect 1494 988 1498 992
rect 901 953 905 957
rect 929 953 933 957
rect 1021 961 1025 965
rect 978 953 982 957
rect 1006 953 1010 957
rect 1046 962 1050 966
rect 1056 962 1060 966
rect 1131 962 1135 966
rect 1056 945 1060 949
rect 1148 945 1152 949
rect 711 932 715 936
rect 790 932 794 936
rect -33 841 -29 845
rect -6 831 -2 835
rect 18 838 22 842
rect 44 845 48 849
rect 68 852 72 856
rect 133 845 137 849
rect 504 845 508 849
rect 131 838 135 842
rect 873 838 877 842
rect 129 831 133 835
rect 1291 831 1295 835
rect 431 754 435 758
rect -322 578 -318 582
rect -476 478 -472 482
rect -630 373 -626 377
rect -784 313 -780 317
rect -707 298 -703 302
rect -769 221 -765 225
rect -692 221 -688 225
rect -553 354 -549 358
rect -615 221 -611 225
rect -538 221 -534 225
rect -399 464 -395 468
rect -461 221 -457 225
rect -384 221 -380 225
rect -245 539 -241 543
rect -307 221 -303 225
rect -230 221 -226 225
rect -169 223 -165 227
rect 136 240 140 244
rect -746 179 -742 183
rect -728 181 -724 185
rect -669 179 -665 183
rect -651 181 -647 185
rect -592 179 -588 183
rect -574 181 -570 185
rect -515 179 -511 183
rect -497 181 -493 185
rect -438 179 -434 183
rect -420 181 -416 185
rect -361 179 -357 183
rect -343 181 -339 185
rect -284 179 -280 183
rect -266 181 -262 185
rect -207 179 -203 183
rect -189 181 -185 185
rect -67 164 -63 168
rect 153 240 157 244
rect 181 240 185 244
rect 34 126 38 130
rect 129 232 133 236
rect 138 232 142 236
rect -67 80 -63 84
rect 230 242 234 246
rect 306 298 310 302
rect 234 208 238 212
rect 61 166 65 170
rect 155 164 159 168
rect 183 164 187 168
rect 140 156 144 160
rect 448 753 452 757
rect 775 754 779 758
rect 710 338 714 342
rect 230 166 234 170
rect 329 164 333 168
rect 476 218 480 222
rect 349 166 353 170
rect 441 206 445 210
rect 499 164 503 168
rect 792 753 796 757
rect 1133 753 1137 757
rect 1106 442 1110 446
rect 519 166 523 170
rect 800 206 804 210
rect 887 164 891 168
rect 1034 215 1038 219
rect 907 166 911 170
rect 999 206 1003 210
rect 1057 164 1061 168
rect 1150 753 1154 757
rect 1479 751 1483 755
rect 1496 753 1500 757
rect 1893 537 1897 541
rect 1077 166 1081 170
rect 1305 206 1309 210
rect 1392 164 1396 168
rect 1539 215 1543 219
rect 1412 166 1416 170
rect 1504 206 1508 210
rect 1562 164 1566 168
rect 1582 166 1586 170
rect 1829 206 1833 210
rect 1916 164 1920 168
rect 2063 576 2067 580
rect 1936 166 1940 170
rect 2028 206 2032 210
rect 2086 164 2090 168
rect 2106 166 2110 170
rect 133 96 137 100
rect -571 0 -567 4
rect -555 2 -551 6
rect -494 0 -490 4
rect -478 2 -474 6
rect -417 0 -413 4
rect -401 2 -397 6
rect -340 0 -336 4
rect -324 2 -320 6
rect 42 45 46 49
rect 58 80 62 84
rect 157 88 161 92
rect 185 88 189 92
rect 142 80 146 84
rect 341 94 345 98
rect 287 58 291 62
rect 271 42 275 46
rect 314 50 318 54
rect 548 92 552 96
rect 330 52 334 56
rect 436 50 440 54
rect 907 92 911 96
rect 456 52 460 56
rect 142 12 146 16
rect 58 6 62 10
rect 159 12 163 16
rect 187 12 191 16
rect 144 4 148 8
rect 606 50 610 54
rect 1106 92 1110 96
rect 626 52 630 56
rect 505 -86 509 -82
rect 490 -94 494 -90
rect 395 -125 399 -121
rect 438 -125 442 -121
rect 573 -121 577 -117
rect 423 -133 427 -129
rect 558 -129 562 -125
rect 505 -169 509 -165
rect 490 -177 494 -173
rect 377 -217 381 -213
rect 994 50 998 54
rect 1412 92 1416 96
rect 1014 52 1018 56
rect 1164 50 1168 54
rect 1611 92 1615 96
rect 1184 52 1188 56
rect 1499 50 1503 54
rect 1936 92 1940 96
rect 1519 52 1523 56
rect 1669 50 1673 54
rect 2135 92 2139 96
rect 1689 52 1693 56
rect 636 -123 640 -119
rect 1018 -86 1022 -82
rect 1003 -94 1007 -90
rect 908 -125 912 -121
rect 951 -125 955 -121
rect 1086 -121 1090 -117
rect 908 -133 912 -129
rect 936 -133 940 -129
rect 1071 -129 1075 -125
rect 1018 -169 1022 -165
rect 1003 -177 1007 -173
rect 906 -215 910 -211
rect 772 -270 776 -266
rect 757 -278 761 -274
rect 1007 -270 1011 -266
rect 992 -278 996 -274
rect 636 -307 640 -303
rect 628 -315 632 -311
rect 662 -307 666 -303
rect 705 -309 709 -305
rect 840 -305 844 -301
rect 662 -319 666 -315
rect 690 -317 694 -313
rect 825 -313 829 -309
rect 881 -307 885 -303
rect 772 -353 776 -349
rect 757 -361 761 -357
rect 869 -398 873 -394
rect 714 -443 718 -439
rect 730 -441 734 -437
rect 940 -309 944 -305
rect 1075 -305 1079 -301
rect 895 -319 899 -315
rect 925 -317 929 -313
rect 1060 -313 1064 -309
rect 1122 -307 1126 -303
rect 1007 -353 1011 -349
rect 992 -361 996 -357
rect 895 -394 899 -390
rect 883 -435 887 -431
rect 938 -443 942 -439
rect 966 -443 970 -439
rect 871 -451 875 -447
rect 923 -451 927 -447
rect 1056 -435 1060 -431
rect 1040 -451 1044 -447
rect 1083 -443 1087 -439
rect 1159 -123 1163 -119
rect 2023 50 2027 54
rect 2043 52 2047 56
rect 2193 50 2197 54
rect 2213 52 2217 56
rect 1524 -86 1528 -82
rect 1509 -94 1513 -90
rect 1414 -125 1418 -121
rect 1457 -125 1461 -121
rect 1592 -121 1596 -117
rect 1414 -133 1418 -129
rect 1442 -133 1446 -129
rect 1577 -129 1581 -125
rect 1524 -169 1528 -165
rect 1509 -177 1513 -173
rect 1412 -215 1416 -211
rect 1295 -270 1299 -266
rect 1280 -278 1284 -274
rect 1530 -270 1534 -266
rect 1515 -278 1519 -274
rect 1159 -307 1163 -303
rect 1151 -315 1155 -311
rect 1185 -307 1189 -303
rect 1228 -309 1232 -305
rect 1363 -305 1367 -301
rect 1185 -319 1189 -315
rect 1213 -317 1217 -313
rect 1348 -313 1352 -309
rect 1404 -307 1408 -303
rect 1295 -353 1299 -349
rect 1280 -361 1284 -357
rect 1392 -398 1396 -394
rect 1237 -443 1241 -439
rect 1253 -441 1257 -437
rect 1463 -309 1467 -305
rect 1598 -305 1602 -301
rect 1418 -319 1422 -315
rect 1448 -317 1452 -313
rect 1583 -313 1587 -309
rect 1645 -307 1649 -303
rect 1530 -353 1534 -349
rect 1515 -361 1519 -357
rect 1418 -394 1422 -390
rect 1406 -435 1410 -431
rect 1461 -443 1465 -439
rect 1489 -443 1493 -439
rect 1394 -451 1398 -447
rect 1446 -451 1450 -447
rect 1579 -435 1583 -431
rect 1563 -451 1567 -447
rect 1606 -443 1610 -439
rect 1682 -123 1686 -119
rect 2048 -86 2052 -82
rect 2033 -94 2037 -90
rect 1938 -125 1942 -121
rect 1981 -125 1985 -121
rect 2116 -121 2120 -117
rect 1938 -133 1942 -129
rect 1966 -133 1970 -129
rect 2101 -129 2105 -125
rect 2048 -169 2052 -165
rect 2033 -177 2037 -173
rect 1936 -215 1940 -211
rect 1818 -270 1822 -266
rect 1803 -278 1807 -274
rect 2053 -270 2057 -266
rect 2038 -278 2042 -274
rect 1682 -307 1686 -303
rect 1674 -315 1678 -311
rect 1708 -307 1712 -303
rect 1751 -309 1755 -305
rect 1886 -305 1890 -301
rect 1708 -319 1712 -315
rect 1736 -317 1740 -313
rect 1871 -313 1875 -309
rect 1927 -307 1931 -303
rect 1818 -353 1822 -349
rect 1803 -361 1807 -357
rect 1915 -398 1919 -394
rect 1760 -443 1764 -439
rect 1776 -441 1780 -437
rect 1986 -309 1990 -305
rect 2121 -305 2125 -301
rect 1941 -319 1945 -315
rect 1971 -317 1975 -313
rect 2106 -313 2110 -309
rect 2168 -307 2172 -303
rect 2053 -353 2057 -349
rect 2038 -361 2042 -357
rect 1941 -394 1945 -390
rect 1929 -435 1933 -431
rect 1984 -443 1988 -439
rect 2012 -443 2016 -439
rect 1917 -451 1921 -447
rect 1969 -451 1973 -447
rect 2102 -435 2106 -431
rect 2086 -451 2090 -447
rect 2129 -443 2133 -439
rect 2205 -123 2209 -119
rect 2341 -270 2345 -266
rect 2326 -278 2330 -274
rect 2576 -270 2580 -266
rect 2561 -278 2565 -274
rect 2205 -307 2209 -303
rect 2197 -315 2201 -311
rect 2231 -307 2235 -303
rect 2274 -309 2278 -305
rect 2409 -305 2413 -301
rect 2231 -319 2235 -315
rect 2259 -317 2263 -313
rect 2394 -313 2398 -309
rect 2450 -307 2454 -303
rect 2341 -353 2345 -349
rect 2326 -361 2330 -357
rect 2438 -398 2442 -394
rect 2283 -443 2287 -439
rect 2299 -441 2303 -437
rect 2509 -309 2513 -305
rect 2644 -305 2648 -301
rect 2464 -319 2468 -315
rect 2494 -317 2498 -313
rect 2629 -313 2633 -309
rect 2691 -307 2695 -303
rect 2576 -353 2580 -349
rect 2561 -361 2565 -357
rect 2464 -394 2468 -390
rect 2452 -435 2456 -431
rect 2507 -443 2511 -439
rect 2535 -443 2539 -439
rect 2440 -451 2444 -447
rect 2492 -451 2496 -447
rect 2625 -435 2629 -431
rect 2609 -451 2613 -447
rect 2652 -443 2656 -439
<< ndcontact >>
rect 10 1524 14 1528
rect 24 1524 28 1528
rect 36 1524 40 1528
rect 51 1524 55 1528
rect 61 1524 65 1528
rect 75 1524 79 1528
rect 87 1524 91 1528
rect 101 1524 105 1528
rect 111 1524 115 1528
rect 125 1524 129 1528
rect 899 1339 903 1343
rect 913 1339 917 1343
rect 925 1339 929 1343
rect 955 1339 959 1343
rect 198 1323 202 1327
rect 212 1323 216 1327
rect 224 1323 228 1327
rect 284 1323 288 1327
rect 305 1322 309 1326
rect 319 1322 323 1326
rect 331 1322 335 1326
rect 361 1322 365 1326
rect 373 1322 377 1326
rect 387 1322 391 1326
rect 555 1325 559 1329
rect 569 1325 573 1329
rect 581 1325 585 1329
rect 626 1325 630 1329
rect 651 1324 655 1328
rect 665 1324 669 1328
rect 677 1324 681 1328
rect 707 1324 711 1328
rect 719 1324 723 1328
rect 733 1324 737 1328
rect 976 1339 980 1343
rect 990 1339 994 1343
rect 1002 1339 1006 1343
rect 1032 1339 1036 1343
rect 1044 1339 1048 1343
rect 1058 1339 1062 1343
rect 1306 1295 1310 1299
rect 1320 1295 1324 1299
rect 1332 1295 1336 1299
rect 1362 1295 1366 1299
rect 1374 1295 1378 1299
rect 1388 1295 1392 1299
rect 632 1185 636 1189
rect 662 1185 666 1189
rect 990 1190 994 1194
rect 1020 1190 1024 1194
rect 1336 1193 1340 1197
rect 1366 1193 1370 1197
rect 288 1177 292 1181
rect 318 1177 322 1181
rect 220 1129 224 1133
rect 250 1129 254 1133
rect 355 1133 359 1137
rect 385 1133 389 1137
rect 564 1137 568 1141
rect 594 1137 598 1141
rect 699 1141 703 1145
rect 729 1141 733 1145
rect 922 1142 926 1146
rect 952 1142 956 1146
rect 1057 1146 1061 1150
rect 1087 1146 1091 1150
rect 1268 1145 1272 1149
rect 163 1120 167 1124
rect 177 1120 181 1124
rect -95 1025 -91 1029
rect -81 1025 -77 1029
rect -69 1025 -65 1029
rect -9 1025 -5 1029
rect 507 1128 511 1132
rect 521 1128 525 1132
rect 288 1094 292 1098
rect 865 1133 869 1137
rect 879 1133 883 1137
rect 318 1094 322 1098
rect 632 1102 636 1106
rect 1298 1145 1302 1149
rect 1403 1149 1407 1153
rect 1433 1149 1437 1153
rect 1211 1136 1215 1140
rect 662 1102 666 1106
rect 990 1107 994 1111
rect 1225 1136 1229 1140
rect 1020 1107 1024 1111
rect 1336 1110 1340 1114
rect 1366 1110 1370 1114
rect 1314 1015 1318 1019
rect 1328 1015 1332 1019
rect 1340 1015 1344 1019
rect 1370 1015 1374 1019
rect 1382 1015 1386 1019
rect 1396 1015 1400 1019
rect 891 972 895 976
rect 905 972 909 976
rect 917 972 921 976
rect 947 972 951 976
rect 527 960 531 964
rect 184 952 188 956
rect 198 952 202 956
rect 210 952 214 956
rect 541 960 545 964
rect 553 960 557 964
rect 598 960 602 964
rect 623 959 627 963
rect 270 952 274 956
rect 291 951 295 955
rect 305 951 309 955
rect 317 951 321 955
rect 347 951 351 955
rect 359 951 363 955
rect 373 951 377 955
rect 637 959 641 963
rect 649 959 653 963
rect 679 959 683 963
rect 691 959 695 963
rect 705 959 709 963
rect 968 972 972 976
rect 982 972 986 976
rect 994 972 998 976
rect 1024 972 1028 976
rect 1036 972 1040 976
rect 1050 972 1054 976
rect -43 861 -39 865
rect -29 861 -25 865
rect -17 861 -13 865
rect -2 861 2 865
rect 8 861 12 865
rect 22 861 26 865
rect 34 861 38 865
rect 48 861 52 865
rect 58 861 62 865
rect 72 861 76 865
rect -792 160 -788 164
rect -762 160 -758 164
rect -750 160 -746 164
rect -736 160 -732 164
rect -715 160 -711 164
rect -685 160 -681 164
rect -673 160 -669 164
rect -659 160 -655 164
rect -638 160 -634 164
rect -608 160 -604 164
rect -596 160 -592 164
rect -582 160 -578 164
rect -561 160 -557 164
rect -531 160 -527 164
rect -519 160 -515 164
rect -505 160 -501 164
rect -484 160 -480 164
rect -454 160 -450 164
rect -442 160 -438 164
rect -428 160 -424 164
rect -407 160 -403 164
rect -377 160 -373 164
rect -365 160 -361 164
rect -351 160 -347 164
rect -330 160 -326 164
rect -300 160 -296 164
rect -288 160 -284 164
rect -274 160 -270 164
rect -253 160 -249 164
rect -223 160 -219 164
rect -211 160 -207 164
rect -197 160 -193 164
rect -71 145 -67 149
rect -57 145 -53 149
rect -71 61 -67 65
rect -57 61 -53 65
rect 135 221 139 225
rect 165 221 169 225
rect 177 221 181 225
rect 191 221 195 225
rect 137 145 141 149
rect 167 145 171 149
rect 179 145 183 149
rect 193 145 197 149
rect 283 145 287 149
rect 313 145 317 149
rect 325 145 329 149
rect 339 145 343 149
rect 453 145 457 149
rect 483 145 487 149
rect 495 145 499 149
rect 509 145 513 149
rect 841 145 845 149
rect 871 145 875 149
rect 883 145 887 149
rect 897 145 901 149
rect 1011 145 1015 149
rect 1041 145 1045 149
rect 1053 145 1057 149
rect 1067 145 1071 149
rect 1346 145 1350 149
rect 1376 145 1380 149
rect 1388 145 1392 149
rect 1402 145 1406 149
rect 1516 145 1520 149
rect 1546 145 1550 149
rect 1558 145 1562 149
rect 1572 145 1576 149
rect 1870 145 1874 149
rect 1900 145 1904 149
rect 1912 145 1916 149
rect 1926 145 1930 149
rect 2040 145 2044 149
rect 2070 145 2074 149
rect 2082 145 2086 149
rect 2096 145 2100 149
rect -617 -19 -613 -15
rect -587 -19 -583 -15
rect -575 -19 -571 -15
rect -561 -19 -557 -15
rect -540 -19 -536 -15
rect -510 -19 -506 -15
rect -498 -19 -494 -15
rect -484 -19 -480 -15
rect -463 -19 -459 -15
rect -433 -19 -429 -15
rect -421 -19 -417 -15
rect -407 -19 -403 -15
rect -386 -19 -382 -15
rect -356 -19 -352 -15
rect -344 -19 -340 -15
rect -330 -19 -326 -15
rect 139 69 143 73
rect 169 69 173 73
rect 181 69 185 73
rect 195 69 199 73
rect 268 31 272 35
rect 282 31 286 35
rect 298 31 302 35
rect 310 31 314 35
rect 324 31 328 35
rect 390 31 394 35
rect 420 31 424 35
rect 432 31 436 35
rect 446 31 450 35
rect 560 31 564 35
rect 590 31 594 35
rect 602 31 606 35
rect 616 31 620 35
rect 141 -7 145 -3
rect 171 -7 175 -3
rect 183 -7 187 -3
rect 197 -7 201 -3
rect 487 -105 491 -101
rect 517 -105 521 -101
rect 420 -144 424 -140
rect 450 -144 454 -140
rect 555 -140 559 -136
rect 585 -140 589 -136
rect 487 -188 491 -184
rect 517 -188 521 -184
rect 948 31 952 35
rect 978 31 982 35
rect 990 31 994 35
rect 1004 31 1008 35
rect 1118 31 1122 35
rect 1148 31 1152 35
rect 1160 31 1164 35
rect 1174 31 1178 35
rect 1453 31 1457 35
rect 1483 31 1487 35
rect 1495 31 1499 35
rect 1509 31 1513 35
rect 1623 31 1627 35
rect 1653 31 1657 35
rect 1665 31 1669 35
rect 1679 31 1683 35
rect 1000 -105 1004 -101
rect 1030 -105 1034 -101
rect 933 -144 937 -140
rect 963 -144 967 -140
rect 1068 -140 1072 -136
rect 1098 -140 1102 -136
rect 1000 -188 1004 -184
rect 1030 -188 1034 -184
rect 754 -289 758 -285
rect 784 -289 788 -285
rect 989 -289 993 -285
rect 687 -328 691 -324
rect 717 -328 721 -324
rect 822 -324 826 -320
rect 852 -324 856 -320
rect 754 -372 758 -368
rect 784 -372 788 -368
rect 668 -462 672 -458
rect 698 -462 702 -458
rect 710 -462 714 -458
rect 724 -462 728 -458
rect 1019 -289 1023 -285
rect 922 -328 926 -324
rect 952 -328 956 -324
rect 1057 -324 1061 -320
rect 1087 -324 1091 -320
rect 989 -372 993 -368
rect 1019 -372 1023 -368
rect 920 -462 924 -458
rect 950 -462 954 -458
rect 962 -462 966 -458
rect 976 -462 980 -458
rect 1037 -462 1041 -458
rect 1051 -462 1055 -458
rect 1067 -462 1071 -458
rect 1079 -462 1083 -458
rect 1093 -462 1097 -458
rect 1977 31 1981 35
rect 2007 31 2011 35
rect 2019 31 2023 35
rect 2033 31 2037 35
rect 2147 31 2151 35
rect 2177 31 2181 35
rect 2189 31 2193 35
rect 2203 31 2207 35
rect 1506 -105 1510 -101
rect 1536 -105 1540 -101
rect 1439 -144 1443 -140
rect 1469 -144 1473 -140
rect 1574 -140 1578 -136
rect 1604 -140 1608 -136
rect 1506 -188 1510 -184
rect 1536 -188 1540 -184
rect 1277 -289 1281 -285
rect 1307 -289 1311 -285
rect 1512 -289 1516 -285
rect 1210 -328 1214 -324
rect 1240 -328 1244 -324
rect 1345 -324 1349 -320
rect 1375 -324 1379 -320
rect 1277 -372 1281 -368
rect 1307 -372 1311 -368
rect 1191 -462 1195 -458
rect 1221 -462 1225 -458
rect 1233 -462 1237 -458
rect 1247 -462 1251 -458
rect 1542 -289 1546 -285
rect 1445 -328 1449 -324
rect 1475 -328 1479 -324
rect 1580 -324 1584 -320
rect 1610 -324 1614 -320
rect 1512 -372 1516 -368
rect 1542 -372 1546 -368
rect 1443 -462 1447 -458
rect 1473 -462 1477 -458
rect 1485 -462 1489 -458
rect 1499 -462 1503 -458
rect 1560 -462 1564 -458
rect 1574 -462 1578 -458
rect 1590 -462 1594 -458
rect 1602 -462 1606 -458
rect 1616 -462 1620 -458
rect 2030 -105 2034 -101
rect 2060 -105 2064 -101
rect 1963 -144 1967 -140
rect 1993 -144 1997 -140
rect 2098 -140 2102 -136
rect 2128 -140 2132 -136
rect 2030 -188 2034 -184
rect 2060 -188 2064 -184
rect 1800 -289 1804 -285
rect 1830 -289 1834 -285
rect 2035 -289 2039 -285
rect 1733 -328 1737 -324
rect 1763 -328 1767 -324
rect 1868 -324 1872 -320
rect 1898 -324 1902 -320
rect 1800 -372 1804 -368
rect 1830 -372 1834 -368
rect 1714 -462 1718 -458
rect 1744 -462 1748 -458
rect 1756 -462 1760 -458
rect 1770 -462 1774 -458
rect 2065 -289 2069 -285
rect 1968 -328 1972 -324
rect 1998 -328 2002 -324
rect 2103 -324 2107 -320
rect 2133 -324 2137 -320
rect 2035 -372 2039 -368
rect 2065 -372 2069 -368
rect 1966 -462 1970 -458
rect 1996 -462 2000 -458
rect 2008 -462 2012 -458
rect 2022 -462 2026 -458
rect 2083 -462 2087 -458
rect 2097 -462 2101 -458
rect 2113 -462 2117 -458
rect 2125 -462 2129 -458
rect 2139 -462 2143 -458
rect 2323 -289 2327 -285
rect 2353 -289 2357 -285
rect 2558 -289 2562 -285
rect 2256 -328 2260 -324
rect 2286 -328 2290 -324
rect 2391 -324 2395 -320
rect 2421 -324 2425 -320
rect 2323 -372 2327 -368
rect 2353 -372 2357 -368
rect 2237 -462 2241 -458
rect 2267 -462 2271 -458
rect 2279 -462 2283 -458
rect 2293 -462 2297 -458
rect 2588 -289 2592 -285
rect 2491 -328 2495 -324
rect 2521 -328 2525 -324
rect 2626 -324 2630 -320
rect 2656 -324 2660 -320
rect 2558 -372 2562 -368
rect 2588 -372 2592 -368
rect 2489 -462 2493 -458
rect 2519 -462 2523 -458
rect 2531 -462 2535 -458
rect 2545 -462 2549 -458
rect 2606 -462 2610 -458
rect 2620 -462 2624 -458
rect 2636 -462 2640 -458
rect 2648 -462 2652 -458
rect 2662 -462 2666 -458
<< pdcontact >>
rect 10 1483 14 1487
rect 24 1483 28 1487
rect 36 1483 40 1487
rect 125 1483 129 1487
rect 899 1299 903 1303
rect 913 1299 917 1303
rect 925 1299 929 1303
rect 940 1299 944 1303
rect 955 1299 959 1303
rect 976 1299 980 1303
rect 990 1299 994 1303
rect 1002 1299 1006 1303
rect 1017 1299 1021 1303
rect 1032 1299 1036 1303
rect 1044 1299 1048 1303
rect 1058 1299 1062 1303
rect 198 1282 202 1286
rect 212 1282 216 1286
rect 224 1282 228 1286
rect 239 1282 243 1286
rect 254 1282 258 1286
rect 269 1282 273 1286
rect 284 1282 288 1286
rect 305 1282 309 1286
rect 319 1282 323 1286
rect 331 1282 335 1286
rect 346 1282 350 1286
rect 361 1282 365 1286
rect 373 1282 377 1286
rect 387 1282 391 1286
rect 555 1284 559 1288
rect 569 1284 573 1288
rect 581 1284 585 1288
rect 596 1284 600 1288
rect 611 1284 615 1288
rect 626 1284 630 1288
rect 651 1284 655 1288
rect 665 1284 669 1288
rect 677 1284 681 1288
rect 692 1284 696 1288
rect 707 1284 711 1288
rect 719 1284 723 1288
rect 733 1284 737 1288
rect 1306 1255 1310 1259
rect 1320 1255 1324 1259
rect 1332 1255 1336 1259
rect 1347 1255 1351 1259
rect 1362 1255 1366 1259
rect 1374 1255 1378 1259
rect 1388 1255 1392 1259
rect 632 1145 636 1149
rect 288 1137 292 1141
rect 303 1137 307 1141
rect 318 1137 322 1141
rect 647 1145 651 1149
rect 990 1150 994 1154
rect 662 1145 666 1149
rect 1005 1150 1009 1154
rect 1020 1150 1024 1154
rect 1336 1153 1340 1157
rect 1351 1153 1355 1157
rect 1366 1153 1370 1157
rect 163 1098 167 1102
rect 177 1098 181 1102
rect 220 1089 224 1093
rect 235 1089 239 1093
rect 250 1089 254 1093
rect 507 1106 511 1110
rect 521 1106 525 1110
rect 355 1093 359 1097
rect 370 1093 374 1097
rect 385 1093 389 1097
rect 564 1097 568 1101
rect 579 1097 583 1101
rect 594 1097 598 1101
rect 865 1111 869 1115
rect 879 1111 883 1115
rect 699 1101 703 1105
rect 714 1101 718 1105
rect 729 1101 733 1105
rect 922 1102 926 1106
rect 937 1102 941 1106
rect 952 1102 956 1106
rect 1211 1114 1215 1118
rect 1225 1114 1229 1118
rect 1057 1106 1061 1110
rect 1072 1106 1076 1110
rect 1087 1106 1091 1110
rect 1268 1105 1272 1109
rect 1283 1105 1287 1109
rect 1298 1105 1302 1109
rect 1403 1109 1407 1113
rect 1418 1109 1422 1113
rect 1433 1109 1437 1113
rect 632 1062 636 1066
rect 647 1062 651 1066
rect 662 1062 666 1066
rect 990 1067 994 1071
rect 1005 1067 1009 1071
rect 1020 1067 1024 1071
rect 1336 1070 1340 1074
rect 1351 1070 1355 1074
rect 1366 1070 1370 1074
rect 288 1054 292 1058
rect 303 1054 307 1058
rect 318 1054 322 1058
rect -95 984 -91 988
rect -81 984 -77 988
rect -69 984 -65 988
rect -54 984 -50 988
rect -39 984 -35 988
rect -24 984 -20 988
rect -9 984 -5 988
rect 1314 975 1318 979
rect 1328 975 1332 979
rect 1340 975 1344 979
rect 1355 975 1359 979
rect 1370 975 1374 979
rect 1382 975 1386 979
rect 1396 975 1400 979
rect 891 932 895 936
rect 905 932 909 936
rect 917 932 921 936
rect 932 932 936 936
rect 947 932 951 936
rect 968 932 972 936
rect 982 932 986 936
rect 994 932 998 936
rect 1009 932 1013 936
rect 1024 932 1028 936
rect 1036 932 1040 936
rect 1050 932 1054 936
rect 527 919 531 923
rect 541 919 545 923
rect 553 919 557 923
rect 568 919 572 923
rect 583 919 587 923
rect 598 919 602 923
rect 623 919 627 923
rect 637 919 641 923
rect 649 919 653 923
rect 664 919 668 923
rect 679 919 683 923
rect 691 919 695 923
rect 705 919 709 923
rect 184 911 188 915
rect 198 911 202 915
rect 210 911 214 915
rect 225 911 229 915
rect 240 911 244 915
rect 255 911 259 915
rect 270 911 274 915
rect 291 911 295 915
rect 305 911 309 915
rect 317 911 321 915
rect 332 911 336 915
rect 347 911 351 915
rect 359 911 363 915
rect 373 911 377 915
rect -43 820 -39 824
rect -29 820 -25 824
rect -17 820 -13 824
rect 72 820 76 824
rect 135 261 139 265
rect 150 261 154 265
rect 165 261 169 265
rect 177 261 181 265
rect 191 261 195 265
rect -792 200 -788 204
rect -777 200 -773 204
rect -762 200 -758 204
rect -750 200 -746 204
rect -736 200 -732 204
rect -715 200 -711 204
rect -700 200 -696 204
rect -685 200 -681 204
rect -673 200 -669 204
rect -659 200 -655 204
rect -638 200 -634 204
rect -623 200 -619 204
rect -608 200 -604 204
rect -596 200 -592 204
rect -582 200 -578 204
rect -561 200 -557 204
rect -546 200 -542 204
rect -531 200 -527 204
rect -519 200 -515 204
rect -505 200 -501 204
rect -484 200 -480 204
rect -469 200 -465 204
rect -454 200 -450 204
rect -442 200 -438 204
rect -428 200 -424 204
rect -407 200 -403 204
rect -392 200 -388 204
rect -377 200 -373 204
rect -365 200 -361 204
rect -351 200 -347 204
rect -330 200 -326 204
rect -315 200 -311 204
rect -300 200 -296 204
rect -288 200 -284 204
rect -274 200 -270 204
rect -253 200 -249 204
rect -238 200 -234 204
rect -223 200 -219 204
rect -211 200 -207 204
rect -197 200 -193 204
rect -71 185 -67 189
rect -57 185 -53 189
rect -71 101 -67 105
rect -57 101 -53 105
rect 137 185 141 189
rect 152 185 156 189
rect 167 185 171 189
rect 179 185 183 189
rect 193 185 197 189
rect 283 185 287 189
rect 298 185 302 189
rect 313 185 317 189
rect 325 185 329 189
rect 339 185 343 189
rect 453 185 457 189
rect 468 185 472 189
rect 483 185 487 189
rect 495 185 499 189
rect 509 185 513 189
rect 841 185 845 189
rect 856 185 860 189
rect 871 185 875 189
rect 883 185 887 189
rect 897 185 901 189
rect 1011 185 1015 189
rect 1026 185 1030 189
rect 1041 185 1045 189
rect 1053 185 1057 189
rect 1067 185 1071 189
rect 1346 185 1350 189
rect 1361 185 1365 189
rect 1376 185 1380 189
rect 1388 185 1392 189
rect 1402 185 1406 189
rect 1516 185 1520 189
rect 1531 185 1535 189
rect 1546 185 1550 189
rect 1558 185 1562 189
rect 1572 185 1576 189
rect 1870 185 1874 189
rect 1885 185 1889 189
rect 1900 185 1904 189
rect 1912 185 1916 189
rect 1926 185 1930 189
rect 2040 185 2044 189
rect 2055 185 2059 189
rect 2070 185 2074 189
rect 2082 185 2086 189
rect 2096 185 2100 189
rect 139 109 143 113
rect 154 109 158 113
rect 169 109 173 113
rect 181 109 185 113
rect 195 109 199 113
rect -617 21 -613 25
rect -602 21 -598 25
rect -587 21 -583 25
rect -575 21 -571 25
rect -561 21 -557 25
rect -540 21 -536 25
rect -525 21 -521 25
rect -510 21 -506 25
rect -498 21 -494 25
rect -484 21 -480 25
rect -463 21 -459 25
rect -448 21 -444 25
rect -433 21 -429 25
rect -421 21 -417 25
rect -407 21 -403 25
rect -386 21 -382 25
rect -371 21 -367 25
rect -356 21 -352 25
rect -344 21 -340 25
rect -330 21 -326 25
rect 268 71 272 75
rect 298 71 302 75
rect 310 71 314 75
rect 324 71 328 75
rect 141 33 145 37
rect 156 33 160 37
rect 171 33 175 37
rect 183 33 187 37
rect 390 71 394 75
rect 405 71 409 75
rect 420 71 424 75
rect 432 71 436 75
rect 446 71 450 75
rect 560 71 564 75
rect 575 71 579 75
rect 590 71 594 75
rect 602 71 606 75
rect 616 71 620 75
rect 197 33 201 37
rect 948 71 952 75
rect 963 71 967 75
rect 978 71 982 75
rect 990 71 994 75
rect 1004 71 1008 75
rect 487 -65 491 -61
rect 502 -65 506 -61
rect 517 -65 521 -61
rect 420 -104 424 -100
rect 435 -104 439 -100
rect 450 -104 454 -100
rect 555 -100 559 -96
rect 570 -100 574 -96
rect 585 -100 589 -96
rect 487 -148 491 -144
rect 502 -148 506 -144
rect 517 -148 521 -144
rect 1118 71 1122 75
rect 1133 71 1137 75
rect 1148 71 1152 75
rect 1160 71 1164 75
rect 1174 71 1178 75
rect 1453 71 1457 75
rect 1468 71 1472 75
rect 1483 71 1487 75
rect 1495 71 1499 75
rect 1509 71 1513 75
rect 1623 71 1627 75
rect 1638 71 1642 75
rect 1653 71 1657 75
rect 1665 71 1669 75
rect 1679 71 1683 75
rect 1977 71 1981 75
rect 1992 71 1996 75
rect 2007 71 2011 75
rect 2019 71 2023 75
rect 2033 71 2037 75
rect 1000 -65 1004 -61
rect 1015 -65 1019 -61
rect 1030 -65 1034 -61
rect 933 -104 937 -100
rect 948 -104 952 -100
rect 963 -104 967 -100
rect 1068 -100 1072 -96
rect 1083 -100 1087 -96
rect 1098 -100 1102 -96
rect 1000 -148 1004 -144
rect 1015 -148 1019 -144
rect 1030 -148 1034 -144
rect 754 -249 758 -245
rect 769 -249 773 -245
rect 784 -249 788 -245
rect 989 -249 993 -245
rect 1004 -249 1008 -245
rect 1019 -249 1023 -245
rect 687 -288 691 -284
rect 702 -288 706 -284
rect 717 -288 721 -284
rect 822 -284 826 -280
rect 837 -284 841 -280
rect 852 -284 856 -280
rect 922 -288 926 -284
rect 937 -288 941 -284
rect 952 -288 956 -284
rect 754 -332 758 -328
rect 769 -332 773 -328
rect 784 -332 788 -328
rect 668 -422 672 -418
rect 683 -422 687 -418
rect 698 -422 702 -418
rect 710 -422 714 -418
rect 724 -422 728 -418
rect 1057 -284 1061 -280
rect 1072 -284 1076 -280
rect 1087 -284 1091 -280
rect 989 -332 993 -328
rect 1004 -332 1008 -328
rect 1019 -332 1023 -328
rect 920 -422 924 -418
rect 935 -422 939 -418
rect 950 -422 954 -418
rect 962 -422 966 -418
rect 976 -422 980 -418
rect 1037 -422 1041 -418
rect 1067 -422 1071 -418
rect 1079 -422 1083 -418
rect 1093 -422 1097 -418
rect 2147 71 2151 75
rect 2162 71 2166 75
rect 2177 71 2181 75
rect 2189 71 2193 75
rect 2203 71 2207 75
rect 1506 -65 1510 -61
rect 1521 -65 1525 -61
rect 1536 -65 1540 -61
rect 1439 -104 1443 -100
rect 1454 -104 1458 -100
rect 1469 -104 1473 -100
rect 1574 -100 1578 -96
rect 1589 -100 1593 -96
rect 1604 -100 1608 -96
rect 1506 -148 1510 -144
rect 1521 -148 1525 -144
rect 1536 -148 1540 -144
rect 1277 -249 1281 -245
rect 1292 -249 1296 -245
rect 1307 -249 1311 -245
rect 1512 -249 1516 -245
rect 1527 -249 1531 -245
rect 1542 -249 1546 -245
rect 1210 -288 1214 -284
rect 1225 -288 1229 -284
rect 1240 -288 1244 -284
rect 1345 -284 1349 -280
rect 1360 -284 1364 -280
rect 1375 -284 1379 -280
rect 1445 -288 1449 -284
rect 1460 -288 1464 -284
rect 1475 -288 1479 -284
rect 1277 -332 1281 -328
rect 1292 -332 1296 -328
rect 1307 -332 1311 -328
rect 1191 -422 1195 -418
rect 1206 -422 1210 -418
rect 1221 -422 1225 -418
rect 1233 -422 1237 -418
rect 1247 -422 1251 -418
rect 1580 -284 1584 -280
rect 1595 -284 1599 -280
rect 1610 -284 1614 -280
rect 1512 -332 1516 -328
rect 1527 -332 1531 -328
rect 1542 -332 1546 -328
rect 1443 -422 1447 -418
rect 1458 -422 1462 -418
rect 1473 -422 1477 -418
rect 1485 -422 1489 -418
rect 1499 -422 1503 -418
rect 1560 -422 1564 -418
rect 1590 -422 1594 -418
rect 1602 -422 1606 -418
rect 1616 -422 1620 -418
rect 2030 -65 2034 -61
rect 2045 -65 2049 -61
rect 2060 -65 2064 -61
rect 1963 -104 1967 -100
rect 1978 -104 1982 -100
rect 1993 -104 1997 -100
rect 2098 -100 2102 -96
rect 2113 -100 2117 -96
rect 2128 -100 2132 -96
rect 2030 -148 2034 -144
rect 2045 -148 2049 -144
rect 2060 -148 2064 -144
rect 1800 -249 1804 -245
rect 1815 -249 1819 -245
rect 1830 -249 1834 -245
rect 2035 -249 2039 -245
rect 2050 -249 2054 -245
rect 2065 -249 2069 -245
rect 1733 -288 1737 -284
rect 1748 -288 1752 -284
rect 1763 -288 1767 -284
rect 1868 -284 1872 -280
rect 1883 -284 1887 -280
rect 1898 -284 1902 -280
rect 1968 -288 1972 -284
rect 1983 -288 1987 -284
rect 1998 -288 2002 -284
rect 1800 -332 1804 -328
rect 1815 -332 1819 -328
rect 1830 -332 1834 -328
rect 1714 -422 1718 -418
rect 1729 -422 1733 -418
rect 1744 -422 1748 -418
rect 1756 -422 1760 -418
rect 1770 -422 1774 -418
rect 2103 -284 2107 -280
rect 2118 -284 2122 -280
rect 2133 -284 2137 -280
rect 2035 -332 2039 -328
rect 2050 -332 2054 -328
rect 2065 -332 2069 -328
rect 1966 -422 1970 -418
rect 1981 -422 1985 -418
rect 1996 -422 2000 -418
rect 2008 -422 2012 -418
rect 2022 -422 2026 -418
rect 2083 -422 2087 -418
rect 2113 -422 2117 -418
rect 2125 -422 2129 -418
rect 2139 -422 2143 -418
rect 2323 -249 2327 -245
rect 2338 -249 2342 -245
rect 2353 -249 2357 -245
rect 2558 -249 2562 -245
rect 2573 -249 2577 -245
rect 2588 -249 2592 -245
rect 2256 -288 2260 -284
rect 2271 -288 2275 -284
rect 2286 -288 2290 -284
rect 2391 -284 2395 -280
rect 2406 -284 2410 -280
rect 2421 -284 2425 -280
rect 2491 -288 2495 -284
rect 2506 -288 2510 -284
rect 2521 -288 2525 -284
rect 2323 -332 2327 -328
rect 2338 -332 2342 -328
rect 2353 -332 2357 -328
rect 2237 -422 2241 -418
rect 2252 -422 2256 -418
rect 2267 -422 2271 -418
rect 2279 -422 2283 -418
rect 2293 -422 2297 -418
rect 2626 -284 2630 -280
rect 2641 -284 2645 -280
rect 2656 -284 2660 -280
rect 2558 -332 2562 -328
rect 2573 -332 2577 -328
rect 2588 -332 2592 -328
rect 2489 -422 2493 -418
rect 2504 -422 2508 -418
rect 2519 -422 2523 -418
rect 2531 -422 2535 -418
rect 2545 -422 2549 -418
rect 2606 -422 2610 -418
rect 2636 -422 2640 -418
rect 2648 -422 2652 -418
rect 2662 -422 2666 -418
<< nbccdiffcontact >>
rect 24 1469 28 1473
rect 913 1285 917 1289
rect 990 1285 994 1289
rect 1058 1285 1062 1289
rect 212 1268 216 1272
rect 319 1268 323 1272
rect 387 1268 391 1272
rect 569 1270 573 1274
rect 665 1270 669 1274
rect 733 1270 737 1274
rect 1320 1241 1324 1245
rect 1388 1241 1392 1245
rect 177 1084 181 1088
rect 521 1092 525 1096
rect 879 1097 883 1101
rect 1225 1100 1229 1104
rect -81 970 -77 974
rect 1328 961 1332 965
rect 1396 961 1400 965
rect 905 918 909 922
rect 982 918 986 922
rect 1050 918 1054 922
rect 541 905 545 909
rect 637 905 641 909
rect 705 905 709 909
rect 198 897 202 901
rect 305 897 309 901
rect 373 897 377 901
rect -29 806 -25 810
rect -750 214 -746 218
rect -673 214 -669 218
rect -596 214 -592 218
rect -519 214 -515 218
rect -442 214 -438 218
rect -365 214 -361 218
rect -288 214 -284 218
rect 177 275 181 279
rect -211 214 -207 218
rect -71 199 -67 203
rect -575 35 -571 39
rect -498 35 -494 39
rect -421 35 -417 39
rect -71 115 -67 119
rect 179 199 183 203
rect 325 199 329 203
rect 495 199 499 203
rect 883 199 887 203
rect 1053 199 1057 203
rect 1388 199 1392 203
rect 1558 199 1562 203
rect 1912 199 1916 203
rect 2082 199 2086 203
rect 181 123 185 127
rect -344 35 -340 39
rect 310 85 314 89
rect 183 47 187 51
rect 432 85 436 89
rect 602 85 606 89
rect 990 85 994 89
rect 1160 85 1164 89
rect 1495 85 1499 89
rect 1665 85 1669 89
rect 2019 85 2023 89
rect 710 -408 714 -404
rect 962 -408 966 -404
rect 1079 -408 1083 -404
rect 2189 85 2193 89
rect 1233 -408 1237 -404
rect 1485 -408 1489 -404
rect 1602 -408 1606 -404
rect 1756 -408 1760 -404
rect 2008 -408 2012 -404
rect 2125 -408 2129 -404
rect 2279 -408 2283 -404
rect 2531 -408 2535 -404
rect 2648 -408 2652 -404
<< m2contact >>
rect 131 1536 135 1540
rect 192 1335 196 1339
rect 393 1334 397 1338
rect 363 1295 367 1299
rect 384 1295 388 1299
rect 395 1268 400 1272
rect 284 1189 288 1193
rect 322 1189 326 1193
rect 216 1141 220 1145
rect 254 1141 258 1145
rect 282 1123 286 1127
rect 323 1123 327 1127
rect 350 1145 354 1149
rect 284 1106 288 1110
rect 352 1079 356 1083
rect 256 1075 260 1079
rect -101 1037 -97 1041
rect -3 1037 1 1041
rect -3 970 1 974
rect 324 1040 328 1044
rect 178 964 182 968
rect 379 963 383 967
rect -49 873 -45 877
rect 349 924 353 928
rect 370 924 374 928
rect 178 897 182 901
rect 379 897 383 901
rect 548 1337 552 1341
rect 739 1336 743 1340
rect 709 1297 713 1301
rect 730 1297 734 1301
rect 547 1270 551 1274
rect 740 1270 744 1274
rect 628 1197 632 1201
rect 666 1197 670 1201
rect 560 1149 564 1153
rect 598 1149 602 1153
rect 626 1131 630 1135
rect 667 1131 671 1135
rect 694 1153 698 1157
rect 628 1114 632 1118
rect 696 1087 700 1091
rect 600 1083 604 1087
rect 626 1048 630 1052
rect 668 1048 672 1052
rect 521 972 525 976
rect 711 971 715 975
rect 681 932 685 936
rect 702 932 706 936
rect 521 905 525 909
rect 712 905 716 909
rect 891 1351 895 1355
rect 1064 1351 1068 1355
rect 1034 1312 1038 1316
rect 1055 1312 1059 1316
rect 894 1285 898 1289
rect 1065 1285 1069 1289
rect 986 1202 990 1206
rect 1024 1202 1028 1206
rect 918 1154 922 1158
rect 956 1154 960 1158
rect 984 1136 988 1140
rect 1025 1136 1029 1140
rect 1052 1158 1056 1162
rect 986 1119 990 1123
rect 1054 1092 1058 1096
rect 958 1088 962 1092
rect 984 1053 988 1057
rect 1026 1053 1030 1057
rect 881 984 885 988
rect 1056 984 1060 988
rect 1026 945 1030 949
rect 1047 945 1051 949
rect 885 918 889 922
rect 1057 918 1061 922
rect 1300 1307 1304 1311
rect 1364 1268 1368 1272
rect 1385 1268 1389 1272
rect 1300 1241 1304 1245
rect 1332 1205 1336 1209
rect 1370 1205 1374 1209
rect 1264 1157 1268 1161
rect 1302 1157 1306 1161
rect 1330 1139 1334 1143
rect 1371 1139 1375 1143
rect 1398 1161 1402 1165
rect 1332 1122 1336 1126
rect 1400 1095 1404 1099
rect 1304 1091 1308 1095
rect 1330 1056 1334 1060
rect 1372 1056 1376 1060
rect 1308 1027 1312 1031
rect 1372 988 1376 992
rect 1393 988 1397 992
rect 1308 961 1312 965
rect 78 806 82 810
rect 27 775 31 779
rect -45 287 -41 291
rect 111 287 115 291
rect 129 275 133 279
rect 197 209 201 213
rect -51 199 -47 203
rect 131 199 135 203
rect -800 148 -796 152
rect -172 148 -168 152
rect -76 133 -72 137
rect -51 115 -47 119
rect 199 133 203 137
rect 230 133 234 137
rect 133 123 137 127
rect -76 49 -72 53
rect 201 57 205 61
rect 135 47 139 51
rect 264 19 268 23
rect 203 -19 207 -15
rect -622 -31 -618 -27
rect -82 -28 -78 -24
rect 216 -28 220 -24
rect 225 -30 229 -26
rect 455 -53 459 -49
rect 968 -53 972 -49
rect 1474 -53 1478 -49
rect 1998 -53 2002 -49
rect 453 -90 457 -86
rect 521 -117 525 -113
rect 455 -156 459 -152
rect 482 -134 486 -130
rect 966 -90 970 -86
rect 1034 -117 1038 -113
rect 551 -152 555 -148
rect 968 -156 972 -152
rect 995 -134 999 -130
rect 1472 -90 1476 -86
rect 1540 -117 1544 -113
rect 1064 -152 1068 -148
rect 1474 -156 1478 -152
rect 1501 -134 1505 -130
rect 1996 -90 2000 -86
rect 2064 -117 2068 -113
rect 1570 -152 1574 -148
rect 1998 -156 2002 -152
rect 2025 -134 2029 -130
rect 2094 -152 2098 -148
rect 465 -198 469 -194
rect 525 -198 529 -194
rect 549 -198 553 -194
rect 978 -198 982 -194
rect 590 -202 594 -198
rect 1038 -198 1042 -194
rect 1062 -198 1066 -194
rect 1484 -198 1488 -194
rect 1544 -198 1548 -194
rect 1568 -198 1572 -194
rect 2008 -198 2012 -194
rect 2068 -198 2072 -194
rect 2092 -198 2096 -194
rect 722 -237 726 -233
rect 957 -237 961 -233
rect 1113 -237 1117 -233
rect 1245 -237 1249 -233
rect 1480 -237 1484 -233
rect 1636 -237 1640 -233
rect 1768 -237 1772 -233
rect 2003 -237 2007 -233
rect 2159 -237 2163 -233
rect 2291 -237 2295 -233
rect 2526 -237 2530 -233
rect 2682 -237 2686 -233
rect 720 -274 724 -270
rect 788 -301 792 -297
rect 955 -274 959 -270
rect 722 -340 726 -336
rect 749 -318 753 -314
rect 1023 -301 1027 -297
rect 818 -336 822 -332
rect 957 -340 961 -336
rect 984 -318 988 -314
rect 1243 -274 1247 -270
rect 1311 -301 1315 -297
rect 1478 -274 1482 -270
rect 1053 -336 1057 -332
rect 1245 -340 1249 -336
rect 1272 -318 1276 -314
rect 1546 -301 1550 -297
rect 1341 -336 1345 -332
rect 1480 -340 1484 -336
rect 1507 -318 1511 -314
rect 1766 -274 1770 -270
rect 1834 -301 1838 -297
rect 2001 -274 2005 -270
rect 1576 -336 1580 -332
rect 1768 -340 1772 -336
rect 1795 -318 1799 -314
rect 2069 -301 2073 -297
rect 1864 -336 1868 -332
rect 2003 -340 2007 -336
rect 2030 -318 2034 -314
rect 2289 -274 2293 -270
rect 2357 -301 2361 -297
rect 2524 -274 2528 -270
rect 2099 -336 2103 -332
rect 2291 -340 2295 -336
rect 2318 -318 2322 -314
rect 2592 -301 2596 -297
rect 2387 -336 2391 -332
rect 2526 -340 2530 -336
rect 2553 -318 2557 -314
rect 2622 -336 2626 -332
rect 732 -382 736 -378
rect 792 -382 796 -378
rect 816 -382 820 -378
rect 967 -382 971 -378
rect 1027 -382 1031 -378
rect 1051 -382 1055 -378
rect 1105 -386 1109 -382
rect 1255 -382 1259 -378
rect 1315 -382 1319 -378
rect 1339 -382 1343 -378
rect 1490 -382 1494 -378
rect 1550 -382 1554 -378
rect 1574 -382 1578 -378
rect 1628 -386 1632 -382
rect 1778 -382 1782 -378
rect 1838 -382 1842 -378
rect 1862 -382 1866 -378
rect 2013 -382 2017 -378
rect 2073 -382 2077 -378
rect 2097 -382 2101 -378
rect 2151 -386 2155 -382
rect 2301 -382 2305 -378
rect 2361 -382 2365 -378
rect 2385 -382 2389 -378
rect 2536 -382 2540 -378
rect 2596 -382 2600 -378
rect 2620 -382 2624 -378
rect 2674 -386 2678 -382
rect 1113 -406 1117 -402
rect 1636 -406 1640 -402
rect 2159 -406 2163 -402
rect 2682 -406 2686 -402
rect 614 -472 618 -468
rect 1105 -472 1109 -468
rect 1628 -472 1632 -468
rect 2151 -472 2155 -468
rect 2674 -472 2678 -468
<< psubstratepcontact >>
rect 9 1536 13 1540
rect 24 1536 28 1540
rect 40 1536 44 1540
rect 70 1536 74 1540
rect 96 1536 100 1540
rect 120 1536 124 1540
rect 197 1335 201 1339
rect 212 1335 216 1339
rect 228 1335 232 1339
rect 279 1335 283 1339
rect 304 1334 308 1338
rect 319 1334 323 1338
rect 335 1334 339 1338
rect 356 1334 360 1338
rect 372 1334 376 1338
rect 387 1334 391 1338
rect 554 1337 558 1341
rect 569 1337 573 1341
rect 585 1337 589 1341
rect 898 1351 902 1355
rect 913 1351 917 1355
rect 929 1351 933 1355
rect 950 1351 954 1355
rect 621 1337 625 1341
rect 650 1336 654 1340
rect 665 1336 669 1340
rect 681 1336 685 1340
rect 702 1336 706 1340
rect 718 1336 722 1340
rect 733 1336 737 1340
rect 975 1351 979 1355
rect 990 1351 994 1355
rect 1006 1351 1010 1355
rect 1027 1351 1031 1355
rect 1043 1351 1047 1355
rect 1058 1351 1062 1355
rect 1305 1307 1309 1311
rect 1320 1307 1324 1311
rect 1336 1307 1340 1311
rect 1357 1307 1361 1311
rect 1373 1307 1377 1311
rect 1388 1307 1392 1311
rect 994 1202 998 1206
rect 1015 1202 1019 1206
rect 1340 1205 1344 1209
rect 1361 1205 1365 1209
rect 636 1197 640 1201
rect 657 1197 661 1201
rect 292 1189 296 1193
rect 313 1189 317 1193
rect 224 1141 228 1145
rect 245 1141 249 1145
rect 568 1149 572 1153
rect 589 1149 593 1153
rect 703 1153 707 1157
rect 724 1153 728 1157
rect 926 1154 930 1158
rect 947 1154 951 1158
rect 1061 1158 1065 1162
rect 1082 1158 1086 1162
rect 1272 1157 1276 1161
rect 1293 1157 1297 1161
rect 1407 1161 1411 1165
rect 1428 1161 1432 1165
rect 359 1145 363 1149
rect 380 1145 384 1149
rect 162 1132 166 1136
rect 177 1132 181 1136
rect 506 1140 510 1144
rect 521 1140 525 1144
rect 864 1145 868 1149
rect 879 1145 883 1149
rect 1210 1148 1214 1152
rect 1225 1148 1229 1152
rect -96 1037 -92 1041
rect -81 1037 -77 1041
rect -65 1037 -61 1041
rect -14 1037 -10 1041
rect 292 1106 296 1110
rect 313 1106 317 1110
rect 636 1114 640 1118
rect 657 1114 661 1118
rect 994 1119 998 1123
rect 1015 1119 1019 1123
rect 1340 1122 1344 1126
rect 1361 1122 1365 1126
rect 1313 1027 1317 1031
rect 1328 1027 1332 1031
rect 1344 1027 1348 1031
rect 1365 1027 1369 1031
rect 1381 1027 1385 1031
rect 1396 1027 1400 1031
rect 183 964 187 968
rect 198 964 202 968
rect 214 964 218 968
rect 526 972 530 976
rect 541 972 545 976
rect 557 972 561 976
rect 265 964 269 968
rect 290 963 294 967
rect 305 963 309 967
rect 321 963 325 967
rect 342 963 346 967
rect 358 963 362 967
rect 373 963 377 967
rect 890 984 894 988
rect 905 984 909 988
rect 921 984 925 988
rect 942 984 946 988
rect 593 972 597 976
rect 622 971 626 975
rect 637 971 641 975
rect 653 971 657 975
rect 674 971 678 975
rect 690 971 694 975
rect 705 971 709 975
rect 967 984 971 988
rect 982 984 986 988
rect 998 984 1002 988
rect 1019 984 1023 988
rect 1035 984 1039 988
rect 1050 984 1054 988
rect -44 873 -40 877
rect -29 873 -25 877
rect -13 873 -9 877
rect 17 873 21 877
rect 43 873 47 877
rect 67 873 71 877
rect -787 148 -783 152
rect -766 148 -762 152
rect -750 148 -746 152
rect -735 148 -731 152
rect -710 148 -706 152
rect -689 148 -685 152
rect -673 148 -669 152
rect -658 148 -654 152
rect -633 148 -629 152
rect -612 148 -608 152
rect -596 148 -592 152
rect -581 148 -577 152
rect -556 148 -552 152
rect -535 148 -531 152
rect -519 148 -515 152
rect -504 148 -500 152
rect -479 148 -475 152
rect -458 148 -454 152
rect -442 148 -438 152
rect -427 148 -423 152
rect -402 148 -398 152
rect -381 148 -377 152
rect -365 148 -361 152
rect -350 148 -346 152
rect -325 148 -321 152
rect -304 148 -300 152
rect -288 148 -284 152
rect -273 148 -269 152
rect -248 148 -244 152
rect -227 148 -223 152
rect -211 148 -207 152
rect -196 148 -192 152
rect -71 133 -67 137
rect -56 133 -52 137
rect 140 209 144 213
rect 161 209 165 213
rect 177 209 181 213
rect 192 209 196 213
rect 142 133 146 137
rect 163 133 167 137
rect 179 133 183 137
rect 194 133 198 137
rect 284 133 288 137
rect 312 133 316 137
rect 325 133 329 137
rect 340 133 344 137
rect 454 133 458 137
rect -71 49 -67 53
rect -56 49 -52 53
rect -612 -31 -608 -27
rect -591 -31 -587 -27
rect -575 -31 -571 -27
rect -560 -31 -556 -27
rect -535 -31 -531 -27
rect -514 -31 -510 -27
rect -498 -31 -494 -27
rect -483 -31 -479 -27
rect -458 -31 -454 -27
rect -437 -31 -433 -27
rect -421 -31 -417 -27
rect -406 -31 -402 -27
rect -381 -31 -377 -27
rect -360 -31 -356 -27
rect -344 -31 -340 -27
rect -329 -31 -325 -27
rect 144 57 148 61
rect 165 57 169 61
rect 181 57 185 61
rect 196 57 200 61
rect 482 133 486 137
rect 495 133 499 137
rect 510 133 514 137
rect 842 133 846 137
rect 870 133 874 137
rect 883 133 887 137
rect 898 133 902 137
rect 1012 133 1016 137
rect 273 19 277 23
rect 294 19 298 23
rect 310 19 314 23
rect 325 19 329 23
rect 391 19 395 23
rect 419 19 423 23
rect 432 19 436 23
rect 447 19 451 23
rect 1040 133 1044 137
rect 1053 133 1057 137
rect 1068 133 1072 137
rect 1347 133 1351 137
rect 1375 133 1379 137
rect 1388 133 1392 137
rect 1403 133 1407 137
rect 1517 133 1521 137
rect 1545 133 1549 137
rect 1558 133 1562 137
rect 1573 133 1577 137
rect 1871 133 1875 137
rect 1899 133 1903 137
rect 1912 133 1916 137
rect 1927 133 1931 137
rect 2041 133 2045 137
rect 561 19 565 23
rect 589 19 593 23
rect 602 19 606 23
rect 617 19 621 23
rect 146 -19 150 -15
rect 167 -19 171 -15
rect 183 -19 187 -15
rect 198 -19 202 -15
rect 492 -117 496 -113
rect 513 -117 517 -113
rect 425 -156 429 -152
rect 446 -156 450 -152
rect 560 -152 564 -148
rect 581 -152 585 -148
rect 492 -200 496 -196
rect 513 -200 517 -196
rect 949 19 953 23
rect 977 19 981 23
rect 990 19 994 23
rect 1005 19 1009 23
rect 1119 19 1123 23
rect 1147 19 1151 23
rect 1160 19 1164 23
rect 1175 19 1179 23
rect 1454 19 1458 23
rect 1482 19 1486 23
rect 1495 19 1499 23
rect 1510 19 1514 23
rect 2069 133 2073 137
rect 2082 133 2086 137
rect 2097 133 2101 137
rect 1624 19 1628 23
rect 1652 19 1656 23
rect 1665 19 1669 23
rect 1680 19 1684 23
rect 1005 -117 1009 -113
rect 1026 -117 1030 -113
rect 938 -156 942 -152
rect 959 -156 963 -152
rect 1073 -152 1077 -148
rect 1094 -152 1098 -148
rect 1005 -200 1009 -196
rect 1026 -200 1030 -196
rect 759 -301 763 -297
rect 780 -301 784 -297
rect 692 -340 696 -336
rect 713 -340 717 -336
rect 827 -336 831 -332
rect 848 -336 852 -332
rect 759 -384 763 -380
rect 780 -384 784 -380
rect 673 -474 677 -470
rect 694 -474 698 -470
rect 710 -474 714 -470
rect 725 -474 729 -470
rect 994 -301 998 -297
rect 1015 -301 1019 -297
rect 927 -340 931 -336
rect 948 -340 952 -336
rect 1062 -336 1066 -332
rect 1083 -336 1087 -332
rect 994 -384 998 -380
rect 1015 -384 1019 -380
rect 925 -474 929 -470
rect 946 -474 950 -470
rect 962 -474 966 -470
rect 977 -474 981 -470
rect 1042 -474 1046 -470
rect 1063 -474 1067 -470
rect 1079 -474 1083 -470
rect 1094 -474 1098 -470
rect 1978 19 1982 23
rect 2006 19 2010 23
rect 2019 19 2023 23
rect 2034 19 2038 23
rect 2148 19 2152 23
rect 2176 19 2180 23
rect 2189 19 2193 23
rect 2204 19 2208 23
rect 1511 -117 1515 -113
rect 1532 -117 1536 -113
rect 1444 -156 1448 -152
rect 1465 -156 1469 -152
rect 1579 -152 1583 -148
rect 1600 -152 1604 -148
rect 1511 -200 1515 -196
rect 1532 -200 1536 -196
rect 1282 -301 1286 -297
rect 1303 -301 1307 -297
rect 1215 -340 1219 -336
rect 1236 -340 1240 -336
rect 1350 -336 1354 -332
rect 1371 -336 1375 -332
rect 1282 -384 1286 -380
rect 1303 -384 1307 -380
rect 1196 -474 1200 -470
rect 1217 -474 1221 -470
rect 1233 -474 1237 -470
rect 1248 -474 1252 -470
rect 1517 -301 1521 -297
rect 1538 -301 1542 -297
rect 1450 -340 1454 -336
rect 1471 -340 1475 -336
rect 1585 -336 1589 -332
rect 1606 -336 1610 -332
rect 1517 -384 1521 -380
rect 1538 -384 1542 -380
rect 1448 -474 1452 -470
rect 1469 -474 1473 -470
rect 1485 -474 1489 -470
rect 1500 -474 1504 -470
rect 1565 -474 1569 -470
rect 1586 -474 1590 -470
rect 1602 -474 1606 -470
rect 1617 -474 1621 -470
rect 2035 -117 2039 -113
rect 2056 -117 2060 -113
rect 1968 -156 1972 -152
rect 1989 -156 1993 -152
rect 2103 -152 2107 -148
rect 2124 -152 2128 -148
rect 2035 -200 2039 -196
rect 2056 -200 2060 -196
rect 1805 -301 1809 -297
rect 1826 -301 1830 -297
rect 1738 -340 1742 -336
rect 1759 -340 1763 -336
rect 1873 -336 1877 -332
rect 1894 -336 1898 -332
rect 1805 -384 1809 -380
rect 1826 -384 1830 -380
rect 1719 -474 1723 -470
rect 1740 -474 1744 -470
rect 1756 -474 1760 -470
rect 1771 -474 1775 -470
rect 2040 -301 2044 -297
rect 2061 -301 2065 -297
rect 1973 -340 1977 -336
rect 1994 -340 1998 -336
rect 2108 -336 2112 -332
rect 2129 -336 2133 -332
rect 2040 -384 2044 -380
rect 2061 -384 2065 -380
rect 1971 -474 1975 -470
rect 1992 -474 1996 -470
rect 2008 -474 2012 -470
rect 2023 -474 2027 -470
rect 2088 -474 2092 -470
rect 2109 -474 2113 -470
rect 2125 -474 2129 -470
rect 2140 -474 2144 -470
rect 2328 -301 2332 -297
rect 2349 -301 2353 -297
rect 2261 -340 2265 -336
rect 2282 -340 2286 -336
rect 2396 -336 2400 -332
rect 2417 -336 2421 -332
rect 2328 -384 2332 -380
rect 2349 -384 2353 -380
rect 2242 -474 2246 -470
rect 2263 -474 2267 -470
rect 2279 -474 2283 -470
rect 2294 -474 2298 -470
rect 2563 -301 2567 -297
rect 2584 -301 2588 -297
rect 2496 -340 2500 -336
rect 2517 -340 2521 -336
rect 2631 -336 2635 -332
rect 2652 -336 2656 -332
rect 2563 -384 2567 -380
rect 2584 -384 2588 -380
rect 2494 -474 2498 -470
rect 2515 -474 2519 -470
rect 2531 -474 2535 -470
rect 2546 -474 2550 -470
rect 2611 -474 2615 -470
rect 2632 -474 2636 -470
rect 2648 -474 2652 -470
rect 2663 -474 2667 -470
<< nsubstratencontact >>
rect 10 1469 14 1473
rect 42 1469 46 1473
rect 70 1469 74 1473
rect 96 1469 100 1473
rect 120 1469 124 1473
rect 899 1285 903 1289
rect 931 1285 935 1289
rect 950 1285 954 1289
rect 976 1285 980 1289
rect 1008 1285 1012 1289
rect 1027 1285 1031 1289
rect 1044 1285 1048 1289
rect 198 1268 202 1272
rect 230 1268 234 1272
rect 279 1268 283 1272
rect 305 1268 309 1272
rect 337 1268 341 1272
rect 356 1268 360 1272
rect 373 1268 377 1272
rect 555 1270 559 1274
rect 587 1270 591 1274
rect 621 1270 625 1274
rect 651 1270 655 1274
rect 683 1270 687 1274
rect 702 1270 706 1274
rect 719 1270 723 1274
rect 1306 1241 1310 1245
rect 1338 1241 1342 1245
rect 1357 1241 1361 1245
rect 1374 1241 1378 1245
rect 294 1123 298 1127
rect 313 1123 317 1127
rect 163 1084 167 1088
rect 638 1131 642 1135
rect 657 1131 661 1135
rect 507 1092 511 1096
rect 996 1136 1000 1140
rect 1015 1136 1019 1140
rect 865 1097 869 1101
rect 1342 1139 1346 1143
rect 1361 1139 1365 1143
rect 1211 1100 1215 1104
rect 570 1083 574 1087
rect 589 1083 593 1087
rect 226 1075 230 1079
rect 245 1075 249 1079
rect 361 1079 365 1083
rect 380 1079 384 1083
rect 705 1087 709 1091
rect 724 1087 728 1091
rect 928 1088 932 1092
rect 947 1088 951 1092
rect 1063 1092 1067 1096
rect 1082 1092 1086 1096
rect 1274 1091 1278 1095
rect 1293 1091 1297 1095
rect 1409 1095 1413 1099
rect 1428 1095 1432 1099
rect 996 1053 1000 1057
rect 1015 1053 1019 1057
rect 1342 1056 1346 1060
rect 1361 1056 1365 1060
rect 638 1048 642 1052
rect 657 1048 661 1052
rect 294 1040 298 1044
rect 313 1040 317 1044
rect -95 970 -91 974
rect -63 970 -59 974
rect -14 970 -10 974
rect 1314 961 1318 965
rect 1346 961 1350 965
rect 1365 961 1369 965
rect 1382 961 1386 965
rect 891 918 895 922
rect 923 918 927 922
rect 942 918 946 922
rect 968 918 972 922
rect 1000 918 1004 922
rect 1019 918 1023 922
rect 1036 918 1040 922
rect 527 905 531 909
rect 559 905 563 909
rect 593 905 597 909
rect 623 905 627 909
rect 655 905 659 909
rect 674 905 678 909
rect 691 905 695 909
rect 184 897 188 901
rect 216 897 220 901
rect 265 897 269 901
rect 291 897 295 901
rect 323 897 327 901
rect 342 897 346 901
rect 359 897 363 901
rect -43 806 -39 810
rect -11 806 -7 810
rect 17 806 21 810
rect 43 806 47 810
rect 67 806 71 810
rect -791 214 -787 218
rect -762 214 -758 218
rect -736 214 -732 218
rect -714 214 -710 218
rect -685 214 -681 218
rect -659 214 -655 218
rect -637 214 -633 218
rect -608 214 -604 218
rect -582 214 -578 218
rect -560 214 -556 218
rect -531 214 -527 218
rect -505 214 -501 218
rect -483 214 -479 218
rect -454 214 -450 218
rect -428 214 -424 218
rect -406 214 -402 218
rect -377 214 -373 218
rect -351 214 -347 218
rect -329 214 -325 218
rect -300 214 -296 218
rect -274 214 -270 218
rect -252 214 -248 218
rect 140 275 144 279
rect 159 275 163 279
rect 191 275 195 279
rect -223 214 -219 218
rect -197 214 -193 218
rect -57 199 -53 203
rect -612 35 -608 39
rect -593 35 -589 39
rect -561 35 -557 39
rect -535 35 -531 39
rect -516 35 -512 39
rect -484 35 -480 39
rect -458 35 -454 39
rect -439 35 -435 39
rect -407 35 -403 39
rect -381 35 -377 39
rect -57 115 -53 119
rect 142 199 146 203
rect 161 199 165 203
rect 193 199 197 203
rect 288 199 292 203
rect 313 199 317 203
rect 339 199 343 203
rect 458 199 462 203
rect 483 199 487 203
rect 509 199 513 203
rect 846 199 850 203
rect 871 199 875 203
rect 897 199 901 203
rect 1016 199 1020 203
rect 1041 199 1045 203
rect 1067 199 1071 203
rect 1351 199 1355 203
rect 1376 199 1380 203
rect 1402 199 1406 203
rect 1521 199 1525 203
rect 1546 199 1550 203
rect 1572 199 1576 203
rect 1875 199 1879 203
rect 1900 199 1904 203
rect 1926 199 1930 203
rect 2045 199 2049 203
rect 2070 199 2074 203
rect 2096 199 2100 203
rect 144 123 148 127
rect 163 123 167 127
rect 195 123 199 127
rect -362 35 -358 39
rect -330 35 -326 39
rect 273 85 277 89
rect 292 85 296 89
rect 324 85 328 89
rect 146 47 150 51
rect 165 47 169 51
rect 197 47 201 51
rect 395 85 399 89
rect 420 85 424 89
rect 446 85 450 89
rect 565 85 569 89
rect 590 85 594 89
rect 616 85 620 89
rect 953 85 957 89
rect 978 85 982 89
rect 1004 85 1008 89
rect 492 -51 496 -47
rect 511 -51 515 -47
rect 425 -90 429 -86
rect 444 -90 448 -86
rect 560 -86 564 -82
rect 579 -86 583 -82
rect 492 -134 496 -130
rect 511 -134 515 -130
rect 1123 85 1127 89
rect 1148 85 1152 89
rect 1174 85 1178 89
rect 1458 85 1462 89
rect 1483 85 1487 89
rect 1509 85 1513 89
rect 1628 85 1632 89
rect 1653 85 1657 89
rect 1679 85 1683 89
rect 1982 85 1986 89
rect 2007 85 2011 89
rect 2033 85 2037 89
rect 1005 -51 1009 -47
rect 1024 -51 1028 -47
rect 938 -90 942 -86
rect 957 -90 961 -86
rect 1073 -86 1077 -82
rect 1092 -86 1096 -82
rect 1005 -134 1009 -130
rect 1024 -134 1028 -130
rect 759 -235 763 -231
rect 778 -235 782 -231
rect 994 -235 998 -231
rect 1013 -235 1017 -231
rect 692 -274 696 -270
rect 711 -274 715 -270
rect 827 -270 831 -266
rect 846 -270 850 -266
rect 927 -274 931 -270
rect 946 -274 950 -270
rect 1062 -270 1066 -266
rect 1081 -270 1085 -266
rect 759 -318 763 -314
rect 778 -318 782 -314
rect 673 -408 677 -404
rect 692 -408 696 -404
rect 724 -408 728 -404
rect 994 -318 998 -314
rect 1013 -318 1017 -314
rect 925 -408 929 -404
rect 944 -408 948 -404
rect 976 -408 980 -404
rect 1042 -408 1046 -404
rect 1061 -408 1065 -404
rect 1093 -408 1097 -404
rect 2152 85 2156 89
rect 2177 85 2181 89
rect 2203 85 2207 89
rect 1511 -51 1515 -47
rect 1530 -51 1534 -47
rect 1444 -90 1448 -86
rect 1463 -90 1467 -86
rect 1579 -86 1583 -82
rect 1598 -86 1602 -82
rect 1511 -134 1515 -130
rect 1530 -134 1534 -130
rect 1282 -235 1286 -231
rect 1301 -235 1305 -231
rect 1517 -235 1521 -231
rect 1536 -235 1540 -231
rect 1215 -274 1219 -270
rect 1234 -274 1238 -270
rect 1350 -270 1354 -266
rect 1369 -270 1373 -266
rect 1450 -274 1454 -270
rect 1469 -274 1473 -270
rect 1585 -270 1589 -266
rect 1604 -270 1608 -266
rect 1282 -318 1286 -314
rect 1301 -318 1305 -314
rect 1196 -408 1200 -404
rect 1215 -408 1219 -404
rect 1247 -408 1251 -404
rect 1517 -318 1521 -314
rect 1536 -318 1540 -314
rect 1448 -408 1452 -404
rect 1467 -408 1471 -404
rect 1499 -408 1503 -404
rect 1565 -408 1569 -404
rect 1584 -408 1588 -404
rect 1616 -408 1620 -404
rect 2035 -51 2039 -47
rect 2054 -51 2058 -47
rect 1968 -90 1972 -86
rect 1987 -90 1991 -86
rect 2103 -86 2107 -82
rect 2122 -86 2126 -82
rect 2035 -134 2039 -130
rect 2054 -134 2058 -130
rect 1805 -235 1809 -231
rect 1824 -235 1828 -231
rect 2040 -235 2044 -231
rect 2059 -235 2063 -231
rect 1738 -274 1742 -270
rect 1757 -274 1761 -270
rect 1873 -270 1877 -266
rect 1892 -270 1896 -266
rect 1973 -274 1977 -270
rect 1992 -274 1996 -270
rect 2108 -270 2112 -266
rect 2127 -270 2131 -266
rect 1805 -318 1809 -314
rect 1824 -318 1828 -314
rect 1719 -408 1723 -404
rect 1738 -408 1742 -404
rect 1770 -408 1774 -404
rect 2040 -318 2044 -314
rect 2059 -318 2063 -314
rect 1971 -408 1975 -404
rect 1990 -408 1994 -404
rect 2022 -408 2026 -404
rect 2088 -408 2092 -404
rect 2107 -408 2111 -404
rect 2139 -408 2143 -404
rect 2328 -235 2332 -231
rect 2347 -235 2351 -231
rect 2563 -235 2567 -231
rect 2582 -235 2586 -231
rect 2261 -274 2265 -270
rect 2280 -274 2284 -270
rect 2396 -270 2400 -266
rect 2415 -270 2419 -266
rect 2496 -274 2500 -270
rect 2515 -274 2519 -270
rect 2631 -270 2635 -266
rect 2650 -270 2654 -266
rect 2328 -318 2332 -314
rect 2347 -318 2351 -314
rect 2242 -408 2246 -404
rect 2261 -408 2265 -404
rect 2293 -408 2297 -404
rect 2563 -318 2567 -314
rect 2582 -318 2586 -314
rect 2494 -408 2498 -404
rect 2513 -408 2517 -404
rect 2545 -408 2549 -404
rect 2611 -408 2615 -404
rect 2630 -408 2634 -404
rect 2662 -408 2666 -404
<< labels >>
rlabel metal1 2704 -439 2704 -439 7 Carry
rlabel polysilicon 2693 -487 2693 -487 1 s3
rlabel polysilicon 2170 -486 2170 -486 1 s2
rlabel polysilicon 1647 -486 1647 -486 1 s1
rlabel polysilicon 1124 -486 1124 -486 1 s0
rlabel metal1 -98 1006 -98 1006 3 E
rlabel metal1 -45 841 -45 841 5 GA
rlabel metal1 8 1504 8 1504 5 GB
rlabel metal1 -63 201 -63 201 1 Vdd
rlabel metal1 -62 51 -62 51 1 gnd
rlabel metal1 -834 302 -834 302 1 b0
rlabel metal1 -817 317 -817 317 1 a0
rlabel metal1 -838 357 -838 357 1 b1
rlabel metal1 -820 377 -820 377 1 a1
rlabel metal1 -839 468 -839 468 3 b2
rlabel metal1 -820 483 -820 483 1 a2
rlabel metal1 -841 543 -841 543 3 b3
rlabel metal1 -818 582 -818 582 1 a3
rlabel metal1 -128 82 -128 82 1 sel0
rlabel metal1 -128 166 -128 166 1 sel1
rlabel polysilicon -551 -43 -551 -43 1 ya0
rlabel polysilicon -474 -43 -474 -43 1 ya1
rlabel polysilicon -397 -43 -397 -43 1 ya2
rlabel polysilicon -320 -43 -320 -43 1 ya3
<< end >>
