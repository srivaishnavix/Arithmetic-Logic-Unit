module New;

initial begin
    $display("Hello, World!");
    $finish; // Finish the simulation
end

endmodule