magic
tech scmos
timestamp 1700583610
<< nwell >>
rect -13 49 100 61
<< polysilicon >>
rect -1 59 2 63
rect 14 59 17 63
rect 29 59 32 63
rect 44 59 47 63
rect 59 59 62 63
rect 86 59 88 63
rect -1 11 2 51
rect 14 11 17 51
rect 29 11 32 51
rect 44 11 47 51
rect 59 11 62 51
rect 86 11 88 51
rect -1 1 2 3
rect 14 1 17 3
rect 29 1 32 3
rect 44 1 47 3
rect 59 1 62 3
rect 86 1 88 3
<< ndiffusion >>
rect -11 9 -1 11
rect -11 5 -9 9
rect -5 5 -1 9
rect -11 3 -1 5
rect 2 3 14 11
rect 17 3 29 11
rect 32 3 44 11
rect 47 3 59 11
rect 62 9 72 11
rect 62 5 66 9
rect 70 5 72 9
rect 62 3 72 5
rect 76 9 86 11
rect 76 5 78 9
rect 82 5 86 9
rect 76 3 86 5
rect 88 9 98 11
rect 88 5 92 9
rect 96 5 98 9
rect 88 3 98 5
<< pdiffusion >>
rect -11 57 -1 59
rect -11 53 -9 57
rect -5 53 -1 57
rect -11 51 -1 53
rect 2 57 14 59
rect 2 53 6 57
rect 10 53 14 57
rect 2 51 14 53
rect 17 57 29 59
rect 17 53 21 57
rect 25 53 29 57
rect 17 51 29 53
rect 32 57 44 59
rect 32 53 36 57
rect 40 53 44 57
rect 32 51 44 53
rect 47 57 59 59
rect 47 53 51 57
rect 55 53 59 57
rect 47 51 59 53
rect 62 57 72 59
rect 62 53 66 57
rect 70 53 72 57
rect 62 51 72 53
rect 76 57 86 59
rect 76 53 78 57
rect 82 53 86 57
rect 76 51 86 53
rect 88 57 98 59
rect 88 53 92 57
rect 96 53 98 57
rect 88 51 98 53
<< metal1 >>
rect -13 67 -4 71
rect 0 67 60 71
rect 64 67 78 71
rect 82 67 92 71
rect 96 67 100 71
rect -9 57 -5 67
rect 66 57 70 67
rect 6 46 10 53
rect 21 46 25 53
rect 36 46 40 53
rect 78 57 82 67
rect 51 46 55 53
rect -15 42 -5 46
rect 6 42 70 46
rect -15 35 10 39
rect -15 28 25 32
rect 66 28 70 42
rect 92 30 96 53
rect -15 21 40 25
rect 66 24 82 28
rect 92 26 100 30
rect -15 14 55 18
rect 66 9 70 24
rect 92 9 96 26
rect -9 -3 -5 5
rect 78 -3 82 5
rect -11 -7 -4 -3
rect 0 -7 62 -3
rect 66 -7 78 -3
rect 82 -7 93 -3
rect 97 -7 100 -3
<< ntransistor >>
rect -1 3 2 11
rect 14 3 17 11
rect 29 3 32 11
rect 44 3 47 11
rect 59 3 62 11
rect 86 3 88 11
<< ptransistor >>
rect -1 51 2 59
rect 14 51 17 59
rect 29 51 32 59
rect 44 51 47 59
rect 59 51 62 59
rect 86 51 88 59
<< polycontact >>
rect -5 42 -1 46
rect 10 35 14 39
rect 25 28 29 32
rect 40 21 44 25
rect 55 14 59 18
rect 82 24 86 28
<< ndcontact >>
rect -9 5 -5 9
rect 66 5 70 9
rect 78 5 82 9
rect 92 5 96 9
<< pdcontact >>
rect -9 53 -5 57
rect 6 53 10 57
rect 21 53 25 57
rect 36 53 40 57
rect 51 53 55 57
rect 66 53 70 57
rect 78 53 82 57
rect 92 53 96 57
<< nbccdiffcontact >>
rect 78 67 82 71
<< psubstratepcontact >>
rect -4 -7 0 -3
rect 62 -7 66 -3
rect 78 -7 82 -3
rect 93 -7 97 -3
<< nsubstratencontact >>
rect -4 67 0 71
rect 60 67 64 71
rect 92 67 96 71
<< labels >>
rlabel metal1 51 69 51 69 5 Vdd
rlabel metal1 -13 44 -13 44 3 Va
rlabel metal1 98 28 98 28 7 Vout
rlabel metal1 53 -5 53 -5 1 gnd
rlabel metal1 -13 37 -13 37 3 Vb
rlabel metal1 -13 30 -13 30 3 Vc
rlabel metal1 -13 23 -13 23 3 Vd
rlabel metal1 -13 16 -13 16 3 Ve
<< end >>
