magic
tech scmos
timestamp 1700582791
<< nwell >>
rect -24 46 74 58
<< polysilicon >>
rect -12 56 -9 60
rect 3 56 6 60
rect 18 56 21 60
rect 33 56 36 60
rect 60 56 62 60
rect -12 15 -9 48
rect 3 15 6 48
rect 18 15 21 48
rect 33 15 36 48
rect 60 15 62 48
rect -12 5 -9 7
rect 3 5 6 7
rect 18 5 21 7
rect 33 5 36 7
rect 60 5 62 7
<< ndiffusion >>
rect -22 13 -12 15
rect -22 9 -20 13
rect -16 9 -12 13
rect -22 7 -12 9
rect -9 7 3 15
rect 6 7 18 15
rect 21 7 33 15
rect 36 13 46 15
rect 36 9 40 13
rect 44 9 46 13
rect 36 7 46 9
rect 50 13 60 15
rect 50 9 52 13
rect 56 9 60 13
rect 50 7 60 9
rect 62 13 72 15
rect 62 9 66 13
rect 70 9 72 13
rect 62 7 72 9
<< pdiffusion >>
rect -22 54 -12 56
rect -22 50 -20 54
rect -16 50 -12 54
rect -22 48 -12 50
rect -9 54 3 56
rect -9 50 -5 54
rect -1 50 3 54
rect -9 48 3 50
rect 6 54 18 56
rect 6 50 10 54
rect 14 50 18 54
rect 6 48 18 50
rect 21 54 33 56
rect 21 50 25 54
rect 29 50 33 54
rect 21 48 33 50
rect 36 54 46 56
rect 36 50 40 54
rect 44 50 46 54
rect 36 48 46 50
rect 50 54 60 56
rect 50 50 52 54
rect 56 50 60 54
rect 50 48 60 50
rect 62 54 72 56
rect 62 50 66 54
rect 70 50 72 54
rect 62 48 72 50
<< metal1 >>
rect -24 64 -15 68
rect -11 64 34 68
rect 38 64 52 68
rect 56 64 66 68
rect 70 64 74 68
rect -20 54 -16 64
rect 40 54 44 64
rect -5 43 -1 50
rect 10 43 14 50
rect 52 54 56 64
rect 25 43 29 50
rect -26 39 -16 43
rect -5 39 44 43
rect -26 32 -1 36
rect 40 32 44 39
rect 66 34 70 50
rect -26 25 14 29
rect 40 28 56 32
rect 66 30 74 34
rect -26 18 29 22
rect 40 13 44 28
rect 66 13 70 30
rect -20 1 -16 9
rect 52 1 56 9
rect -22 -3 -15 1
rect -11 -3 36 1
rect 40 -3 52 1
rect 56 -3 67 1
rect 71 -3 74 1
<< ntransistor >>
rect -12 7 -9 15
rect 3 7 6 15
rect 18 7 21 15
rect 33 7 36 15
rect 60 7 62 15
<< ptransistor >>
rect -12 48 -9 56
rect 3 48 6 56
rect 18 48 21 56
rect 33 48 36 56
rect 60 48 62 56
<< polycontact >>
rect -16 39 -12 43
rect -1 32 3 36
rect 14 25 18 29
rect 29 18 33 22
rect 56 28 60 32
<< ndcontact >>
rect -20 9 -16 13
rect 40 9 44 13
rect 52 9 56 13
rect 66 9 70 13
<< pdcontact >>
rect -20 50 -16 54
rect -5 50 -1 54
rect 10 50 14 54
rect 25 50 29 54
rect 40 50 44 54
rect 52 50 56 54
rect 66 50 70 54
<< nbccdiffcontact >>
rect 52 64 56 68
<< psubstratepcontact >>
rect -15 -3 -11 1
rect 36 -3 40 1
rect 52 -3 56 1
rect 67 -3 71 1
<< nsubstratencontact >>
rect -15 64 -11 68
rect 34 64 38 68
rect 66 64 70 68
<< labels >>
rlabel metal1 -24 41 -24 41 3 Va
rlabel metal1 -24 34 -24 34 3 Vb
rlabel metal1 -24 27 -24 27 3 Vc
rlabel metal1 -24 20 -24 20 3 Vd
rlabel metal1 72 32 72 32 7 Vout
rlabel metal1 25 66 25 66 5 Vdd
rlabel metal1 27 -1 27 -1 1 gnd
<< end >>
