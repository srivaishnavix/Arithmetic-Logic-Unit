FullAdder gate implementation using AND OR gates

.include TSMC_180nm.txt
.include NAND.sub
.include NOT.sub
.include AND.sub
.include OR.sub
.include XOR.sub
.include XNOR.sub
.include FullAdder.sub


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a node_a gnd dc 'supply'
V_in_b node_b gnd dc 'supply'
V_in_c node_c gnd dc    0

X1 node_a node_b node_c node_s node_cout node_x gnd FullAdder

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_a) v(node_b)+2 v(node_c)+4 v(node_s)+6 v(node_cout)+8
.end
.endc