magic
tech scmos
timestamp 1700587889
<< nwell >>
rect -48 55 -6 67
rect -115 16 -73 28
rect 20 20 62 32
rect 93 11 119 23
rect -48 -28 -6 -16
<< polysilicon >>
rect -36 65 -33 69
rect -21 65 -18 69
rect -36 34 -33 57
rect -21 42 -18 57
rect -22 38 -18 42
rect -37 30 -33 34
rect -103 26 -100 30
rect -88 26 -85 30
rect -36 25 -33 30
rect -21 25 -18 38
rect 32 30 35 34
rect 47 30 50 34
rect -103 -5 -100 18
rect -88 3 -85 18
rect -36 15 -33 17
rect -21 15 -18 17
rect -89 -1 -85 3
rect 32 -1 35 22
rect 47 7 50 22
rect 105 21 107 25
rect 46 3 50 7
rect -104 -9 -100 -5
rect -103 -14 -100 -9
rect -88 -14 -85 -1
rect 31 -5 35 -1
rect 32 -10 35 -5
rect 47 -10 50 3
rect 105 -1 107 13
rect -36 -18 -33 -14
rect -21 -18 -18 -14
rect 105 -11 107 -9
rect -103 -24 -100 -22
rect -88 -24 -85 -22
rect 32 -20 35 -18
rect 47 -20 50 -18
rect -36 -49 -33 -26
rect -21 -41 -18 -26
rect -22 -45 -18 -41
rect -37 -53 -33 -49
rect -36 -58 -33 -53
rect -21 -58 -18 -45
rect -36 -68 -33 -66
rect -21 -68 -18 -66
<< ndiffusion >>
rect -46 23 -36 25
rect -46 19 -44 23
rect -40 19 -36 23
rect -46 17 -36 19
rect -33 17 -21 25
rect -18 23 -8 25
rect -18 19 -14 23
rect -10 19 -8 23
rect -18 17 -8 19
rect 95 -3 105 -1
rect 95 -7 97 -3
rect 101 -7 105 -3
rect 95 -9 105 -7
rect 107 -3 117 -1
rect 107 -7 111 -3
rect 115 -7 117 -3
rect 107 -9 117 -7
rect 22 -12 32 -10
rect -113 -16 -103 -14
rect -113 -20 -111 -16
rect -107 -20 -103 -16
rect -113 -22 -103 -20
rect -100 -22 -88 -14
rect -85 -16 -75 -14
rect -85 -20 -81 -16
rect -77 -20 -75 -16
rect 22 -16 24 -12
rect 28 -16 32 -12
rect 22 -18 32 -16
rect 35 -18 47 -10
rect 50 -12 60 -10
rect 50 -16 54 -12
rect 58 -16 60 -12
rect 50 -18 60 -16
rect -85 -22 -75 -20
rect -46 -60 -36 -58
rect -46 -64 -44 -60
rect -40 -64 -36 -60
rect -46 -66 -36 -64
rect -33 -66 -21 -58
rect -18 -60 -8 -58
rect -18 -64 -14 -60
rect -10 -64 -8 -60
rect -18 -66 -8 -64
<< pdiffusion >>
rect -46 63 -36 65
rect -46 59 -44 63
rect -40 59 -36 63
rect -46 57 -36 59
rect -33 63 -21 65
rect -33 59 -29 63
rect -25 59 -21 63
rect -33 57 -21 59
rect -18 63 -8 65
rect -18 59 -14 63
rect -10 59 -8 63
rect -18 57 -8 59
rect -113 24 -103 26
rect -113 20 -111 24
rect -107 20 -103 24
rect -113 18 -103 20
rect -100 24 -88 26
rect -100 20 -96 24
rect -92 20 -88 24
rect -100 18 -88 20
rect -85 24 -75 26
rect 22 28 32 30
rect -85 20 -81 24
rect -77 20 -75 24
rect -85 18 -75 20
rect 22 24 24 28
rect 28 24 32 28
rect 22 22 32 24
rect 35 28 47 30
rect 35 24 39 28
rect 43 24 47 28
rect 35 22 47 24
rect 50 28 60 30
rect 50 24 54 28
rect 58 24 60 28
rect 50 22 60 24
rect 95 19 105 21
rect 95 15 97 19
rect 101 15 105 19
rect 95 13 105 15
rect 107 19 117 21
rect 107 15 111 19
rect 115 15 117 19
rect 107 13 117 15
rect -46 -20 -36 -18
rect -46 -24 -44 -20
rect -40 -24 -36 -20
rect -46 -26 -36 -24
rect -33 -20 -21 -18
rect -33 -24 -29 -20
rect -25 -24 -21 -20
rect -33 -26 -21 -24
rect -18 -20 -8 -18
rect -18 -24 -14 -20
rect -10 -24 -8 -20
rect -18 -26 -8 -24
<< metal1 >>
rect -46 73 -39 77
rect -35 73 -20 77
rect -16 73 -6 77
rect -44 63 -40 73
rect -14 63 -10 73
rect -29 50 -25 59
rect -29 46 -10 50
rect -123 42 -48 46
rect -14 42 -10 46
rect -123 3 -118 42
rect -52 38 -26 42
rect -14 38 6 42
rect 22 38 29 42
rect 33 38 48 42
rect 52 38 93 42
rect -115 34 -106 38
rect -102 34 -87 38
rect -83 34 -78 38
rect -111 24 -107 34
rect -81 24 -77 34
rect -61 30 -41 34
rect -96 11 -92 20
rect -96 7 -77 11
rect -81 3 -77 7
rect -61 3 -57 30
rect -14 23 -10 38
rect -44 11 -40 19
rect -46 7 -39 11
rect -35 7 -18 11
rect -14 7 -10 11
rect 2 7 6 38
rect 24 28 28 38
rect 54 28 58 38
rect 89 33 93 38
rect 89 29 97 33
rect 101 29 111 33
rect 115 29 119 33
rect 39 15 43 24
rect 97 19 101 29
rect 39 11 58 15
rect 54 7 58 11
rect 111 8 115 15
rect 2 3 42 7
rect 54 3 101 7
rect 111 4 123 8
rect -134 -1 -93 3
rect -81 -1 -57 3
rect -134 -9 -108 -5
rect -121 -36 -116 -9
rect -81 -16 -77 -1
rect -111 -28 -107 -20
rect -113 -32 -106 -28
rect -102 -32 -85 -28
rect -81 -32 -76 -28
rect -121 -40 -66 -36
rect -71 -49 -66 -40
rect -61 -41 -57 -1
rect 2 -5 27 -1
rect -45 -10 -39 -6
rect -35 -10 -20 -6
rect -16 -10 -8 -6
rect -44 -20 -40 -10
rect -14 -20 -10 -10
rect -29 -33 -25 -24
rect -29 -37 -10 -33
rect -14 -41 -10 -37
rect 2 -41 6 -5
rect 54 -12 58 3
rect 111 -3 115 4
rect 97 -15 101 -7
rect 24 -24 28 -16
rect 91 -19 97 -15
rect 101 -19 112 -15
rect 116 -19 119 -15
rect 24 -28 29 -24
rect 33 -28 50 -24
rect 54 -32 58 -24
rect 91 -32 95 -19
rect 54 -36 95 -32
rect -61 -45 -26 -41
rect -14 -45 6 -41
rect -71 -53 -41 -49
rect -14 -60 -10 -45
rect -44 -72 -40 -64
rect -44 -76 -39 -72
rect -35 -76 -18 -72
rect -14 -76 -10 -72
rect -29 -80 -25 -76
<< metal2 >>
rect -76 73 -50 77
rect -76 38 -72 73
rect -5 46 70 50
rect -74 34 -64 38
rect -68 -6 -64 34
rect -5 11 -1 46
rect -6 7 -1 11
rect 11 38 18 42
rect 11 -6 15 38
rect -68 -10 -49 -6
rect -4 -10 15 -6
rect 66 -24 70 46
rect 18 -28 20 -24
rect 62 -28 70 -24
rect -72 -32 -62 -28
rect -66 -72 -62 -32
rect 18 -72 22 -28
rect -66 -76 -48 -72
rect -6 -76 22 -72
<< ntransistor >>
rect -36 17 -33 25
rect -21 17 -18 25
rect 105 -9 107 -1
rect -103 -22 -100 -14
rect -88 -22 -85 -14
rect 32 -18 35 -10
rect 47 -18 50 -10
rect -36 -66 -33 -58
rect -21 -66 -18 -58
<< ptransistor >>
rect -36 57 -33 65
rect -21 57 -18 65
rect -103 18 -100 26
rect -88 18 -85 26
rect 32 22 35 30
rect 47 22 50 30
rect 105 13 107 21
rect -36 -26 -33 -18
rect -21 -26 -18 -18
<< polycontact >>
rect -26 38 -22 42
rect -41 30 -37 34
rect -93 -1 -89 3
rect 42 3 46 7
rect 101 3 105 7
rect -108 -9 -104 -5
rect 27 -5 31 -1
rect -26 -45 -22 -41
rect -41 -53 -37 -49
<< ndcontact >>
rect -44 19 -40 23
rect -14 19 -10 23
rect 97 -7 101 -3
rect 111 -7 115 -3
rect -111 -20 -107 -16
rect -81 -20 -77 -16
rect 24 -16 28 -12
rect 54 -16 58 -12
rect -44 -64 -40 -60
rect -14 -64 -10 -60
<< pdcontact >>
rect -44 59 -40 63
rect -29 59 -25 63
rect -14 59 -10 63
rect -111 20 -107 24
rect -96 20 -92 24
rect -81 20 -77 24
rect 24 24 28 28
rect 39 24 43 28
rect 54 24 58 28
rect 97 15 101 19
rect 111 15 115 19
rect -44 -24 -40 -20
rect -29 -24 -25 -20
rect -14 -24 -10 -20
<< nbccdiffcontact >>
rect 97 29 101 33
<< m2contact >>
rect -50 73 -46 77
rect 18 38 22 42
rect -78 34 -74 38
rect -10 7 -6 11
rect -76 -32 -72 -28
rect -49 -10 -45 -6
rect -8 -10 -4 -6
rect 20 -28 24 -24
rect 58 -28 62 -24
rect -48 -76 -44 -72
rect -10 -76 -6 -72
<< psubstratepcontact >>
rect -39 7 -35 11
rect -18 7 -14 11
rect 97 -19 101 -15
rect 112 -19 116 -15
rect -106 -32 -102 -28
rect -85 -32 -81 -28
rect 29 -28 33 -24
rect 50 -28 54 -24
rect -39 -76 -35 -72
rect -18 -76 -14 -72
<< nsubstratencontact >>
rect -39 73 -35 77
rect -20 73 -16 77
rect -106 34 -102 38
rect -87 34 -83 38
rect 29 38 33 42
rect 48 38 52 42
rect 111 29 115 33
rect -39 -10 -35 -6
rect -20 -10 -16 -6
<< end >>
