* SPICE3 file created from 4ANDGAT.ext - technology: scmos

.include TSMC_180nm.txt

.param SUPPLY = 1
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd Vdd gnd 'SUPPLY'

.option scale=1u

M1000 a_n9_48# Vc a_n9_48# w_n24_46# CMOSP w=8 l=3
+  ad=48p pd=20u as=0.288n ps=0.12m
M1001 a_21_7# Vc a_6_7# Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=48p ps=20u
M1002 Vout a_n9_48# Vdd w_n24_46# CMOSP w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1003 a_n9_7# Va gnd Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
M1004 a_6_7# Vb a_n9_7# Gnd CMOSN w=8 l=3
+  ad=48p pd=20u as=48p ps=20u
M1005 Vout a_n9_48# gnd Gnd CMOSN w=8 l=2
+  ad=80p pd=36u as=80p ps=36u
M1006 a_n9_48# Vb a_n9_48# w_n24_46# CMOSP w=8 l=3
+  ad=48p pd=20u as=0 ps=0
M1007 a_n9_48# Vd a_21_7# Gnd CMOSN w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1008 Vdd Vd a_n9_48# w_n24_46# CMOSP w=8 l=3
+  ad=80p pd=36u as=48p ps=20u
M1009 a_n9_48# Va Vdd w_n24_46# CMOSP w=8 l=3
+  ad=48p pd=20u as=80p ps=36u
C0 gnd 0 17.296f 
C1 Vout 0 6.58f 
C2 a_n9_48# 0 27.174f 
C3 Vd 0 21.687f 
C4 Vc 0 19.431f 
C5 Vb 0 17.175001f 
C6 Va 0 14.919f 
C7 Vdd 0 18.8f 


Va Va gnd 1
Vb Vb gnd 1
Vc Vc gnd 0
Vd Vd gnd 1


.tran 1n 800n
.control

run
set color0 = rgb:f/f/e
set color1 = black
plot v(Va) v(Vb)+2 v(Vc)+4 v(Vd)+6 v(Vout)+8 
.end
.endc