magic
tech scmos
timestamp 1701007510
<< nwell >>
rect -30 55 12 67
rect -97 16 -55 28
rect 38 20 80 32
rect -30 -28 12 -16
<< polysilicon >>
rect -18 65 -15 69
rect -3 65 0 69
rect -18 34 -15 57
rect -3 42 0 57
rect -4 38 0 42
rect -19 30 -15 34
rect -85 26 -82 30
rect -70 26 -67 30
rect -18 25 -15 30
rect -3 25 0 38
rect 50 30 53 34
rect 65 30 68 34
rect -85 -5 -82 18
rect -70 3 -67 18
rect -18 15 -15 17
rect -3 15 0 17
rect -71 -1 -67 3
rect 50 -1 53 22
rect 65 7 68 22
rect 64 3 68 7
rect -86 -9 -82 -5
rect -85 -14 -82 -9
rect -70 -14 -67 -1
rect 49 -5 53 -1
rect 50 -10 53 -5
rect 65 -10 68 3
rect -18 -18 -15 -14
rect -3 -18 0 -14
rect -85 -24 -82 -22
rect -70 -24 -67 -22
rect 50 -20 53 -18
rect 65 -20 68 -18
rect -18 -49 -15 -26
rect -3 -41 0 -26
rect -4 -45 0 -41
rect -19 -53 -15 -49
rect -18 -58 -15 -53
rect -3 -58 0 -45
rect -18 -68 -15 -66
rect -3 -68 0 -66
<< ndiffusion >>
rect -28 23 -18 25
rect -28 19 -26 23
rect -22 19 -18 23
rect -28 17 -18 19
rect -15 17 -3 25
rect 0 23 10 25
rect 0 19 4 23
rect 8 19 10 23
rect 0 17 10 19
rect 40 -12 50 -10
rect -95 -16 -85 -14
rect -95 -20 -93 -16
rect -89 -20 -85 -16
rect -95 -22 -85 -20
rect -82 -22 -70 -14
rect -67 -16 -57 -14
rect -67 -20 -63 -16
rect -59 -20 -57 -16
rect 40 -16 42 -12
rect 46 -16 50 -12
rect 40 -18 50 -16
rect 53 -18 65 -10
rect 68 -12 78 -10
rect 68 -16 72 -12
rect 76 -16 78 -12
rect 68 -18 78 -16
rect -67 -22 -57 -20
rect -28 -60 -18 -58
rect -28 -64 -26 -60
rect -22 -64 -18 -60
rect -28 -66 -18 -64
rect -15 -66 -3 -58
rect 0 -60 10 -58
rect 0 -64 4 -60
rect 8 -64 10 -60
rect 0 -66 10 -64
<< pdiffusion >>
rect -28 63 -18 65
rect -28 59 -26 63
rect -22 59 -18 63
rect -28 57 -18 59
rect -15 63 -3 65
rect -15 59 -11 63
rect -7 59 -3 63
rect -15 57 -3 59
rect 0 63 10 65
rect 0 59 4 63
rect 8 59 10 63
rect 0 57 10 59
rect -95 24 -85 26
rect -95 20 -93 24
rect -89 20 -85 24
rect -95 18 -85 20
rect -82 24 -70 26
rect -82 20 -78 24
rect -74 20 -70 24
rect -82 18 -70 20
rect -67 24 -57 26
rect 40 28 50 30
rect -67 20 -63 24
rect -59 20 -57 24
rect -67 18 -57 20
rect 40 24 42 28
rect 46 24 50 28
rect 40 22 50 24
rect 53 28 65 30
rect 53 24 57 28
rect 61 24 65 28
rect 53 22 65 24
rect 68 28 78 30
rect 68 24 72 28
rect 76 24 78 28
rect 68 22 78 24
rect -28 -20 -18 -18
rect -28 -24 -26 -20
rect -22 -24 -18 -20
rect -28 -26 -18 -24
rect -15 -20 -3 -18
rect -15 -24 -11 -20
rect -7 -24 -3 -20
rect -15 -26 -3 -24
rect 0 -20 10 -18
rect 0 -24 4 -20
rect 8 -24 10 -20
rect 0 -26 10 -24
<< metal1 >>
rect -118 75 -21 77
rect -118 73 -58 75
rect -54 73 -21 75
rect -17 73 -2 77
rect 2 73 107 77
rect -26 63 -22 73
rect 4 63 8 73
rect -11 50 -7 59
rect -11 46 8 50
rect -105 42 -30 46
rect 4 42 8 46
rect 59 42 63 73
rect -105 3 -100 42
rect -34 38 -8 42
rect 4 38 24 42
rect 40 38 47 42
rect 51 38 66 42
rect 70 38 80 42
rect -97 34 -88 38
rect -84 34 -69 38
rect -65 34 -60 38
rect -93 24 -89 34
rect -63 24 -59 34
rect -43 30 -23 34
rect -78 11 -74 20
rect -78 7 -59 11
rect -63 3 -59 7
rect -43 3 -39 30
rect 4 23 8 38
rect -26 11 -22 19
rect -28 7 -21 11
rect -17 7 0 11
rect 4 7 8 11
rect 20 7 24 38
rect 42 28 46 38
rect 72 28 76 38
rect 57 15 61 24
rect 57 11 76 15
rect 72 7 76 11
rect 20 3 60 7
rect 72 3 107 7
rect -116 -1 -75 3
rect -63 -1 -39 3
rect -116 -9 -90 -5
rect -103 -36 -98 -9
rect -63 -16 -59 -1
rect -93 -28 -89 -20
rect -95 -32 -88 -28
rect -84 -32 -67 -28
rect -63 -32 -58 -28
rect -103 -40 -48 -36
rect -53 -49 -48 -40
rect -43 -41 -39 -1
rect 20 -5 45 -1
rect -27 -10 -21 -6
rect -17 -10 -2 -6
rect 2 -10 10 -6
rect -26 -20 -22 -10
rect 4 -20 8 -10
rect -11 -33 -7 -24
rect -11 -37 8 -33
rect 4 -41 8 -37
rect 20 -41 24 -5
rect 72 -12 76 3
rect 42 -24 46 -16
rect 42 -28 47 -24
rect 51 -28 68 -24
rect 72 -28 76 -24
rect -43 -45 -8 -41
rect 4 -45 24 -41
rect -53 -53 -23 -49
rect 4 -60 8 -45
rect -118 -74 -48 -72
rect -26 -72 -22 -64
rect -44 -74 -21 -72
rect -118 -76 -21 -74
rect -17 -76 0 -72
rect 4 -74 12 -72
rect 16 -74 36 -72
rect 40 -74 108 -72
rect 4 -76 108 -74
<< metal2 >>
rect -58 38 -54 71
rect -56 34 -46 38
rect -50 -6 -46 34
rect -50 -10 -31 -6
rect -54 -32 -44 -28
rect -48 -70 -44 -32
rect 12 -70 16 11
rect 36 -28 38 -24
rect 36 -70 40 -28
<< ntransistor >>
rect -18 17 -15 25
rect -3 17 0 25
rect -85 -22 -82 -14
rect -70 -22 -67 -14
rect 50 -18 53 -10
rect 65 -18 68 -10
rect -18 -66 -15 -58
rect -3 -66 0 -58
<< ptransistor >>
rect -18 57 -15 65
rect -3 57 0 65
rect -85 18 -82 26
rect -70 18 -67 26
rect 50 22 53 30
rect 65 22 68 30
rect -18 -26 -15 -18
rect -3 -26 0 -18
<< polycontact >>
rect -8 38 -4 42
rect -23 30 -19 34
rect -75 -1 -71 3
rect 60 3 64 7
rect -90 -9 -86 -5
rect 45 -5 49 -1
rect -8 -45 -4 -41
rect -23 -53 -19 -49
<< ndcontact >>
rect -26 19 -22 23
rect 4 19 8 23
rect -93 -20 -89 -16
rect -63 -20 -59 -16
rect 42 -16 46 -12
rect 72 -16 76 -12
rect -26 -64 -22 -60
rect 4 -64 8 -60
<< pdcontact >>
rect -26 59 -22 63
rect -11 59 -7 63
rect 4 59 8 63
rect -93 20 -89 24
rect -78 20 -74 24
rect -63 20 -59 24
rect 42 24 46 28
rect 57 24 61 28
rect 72 24 76 28
rect -26 -24 -22 -20
rect -11 -24 -7 -20
rect 4 -24 8 -20
<< m2contact >>
rect -58 71 -54 75
rect -60 34 -56 38
rect 8 7 12 11
rect -58 -32 -54 -28
rect -31 -10 -27 -6
rect 38 -28 42 -24
rect -48 -74 -44 -70
rect 12 -74 16 -70
rect 36 -74 40 -70
<< psubstratepcontact >>
rect -21 7 -17 11
rect 0 7 4 11
rect -88 -32 -84 -28
rect -67 -32 -63 -28
rect 47 -28 51 -24
rect 68 -28 72 -24
rect -21 -76 -17 -72
rect 0 -76 4 -72
<< nsubstratencontact >>
rect -21 73 -17 77
rect -2 73 2 77
rect -88 34 -84 38
rect -69 34 -65 38
rect 47 38 51 42
rect 66 38 70 42
rect -21 -10 -17 -6
rect -2 -10 2 -6
<< end >>
